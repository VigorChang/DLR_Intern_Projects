-- soc.vhd

-- Generated using ACDS version 15.0 145

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc is
	port (
		clk_clk            : in    std_logic                     := '0';             --    clk.clk
		memory_mem_a       : out   std_logic_vector(14 downto 0);                    -- memory.mem_a
		memory_mem_ba      : out   std_logic_vector(2 downto 0);                     --       .mem_ba
		memory_mem_ck      : out   std_logic;                                        --       .mem_ck
		memory_mem_ck_n    : out   std_logic;                                        --       .mem_ck_n
		memory_mem_cke     : out   std_logic;                                        --       .mem_cke
		memory_mem_cs_n    : out   std_logic;                                        --       .mem_cs_n
		memory_mem_ras_n   : out   std_logic;                                        --       .mem_ras_n
		memory_mem_cas_n   : out   std_logic;                                        --       .mem_cas_n
		memory_mem_we_n    : out   std_logic;                                        --       .mem_we_n
		memory_mem_reset_n : out   std_logic;                                        --       .mem_reset_n
		memory_mem_dq      : inout std_logic_vector(31 downto 0) := (others => '0'); --       .mem_dq
		memory_mem_dqs     : inout std_logic_vector(3 downto 0)  := (others => '0'); --       .mem_dqs
		memory_mem_dqs_n   : inout std_logic_vector(3 downto 0)  := (others => '0'); --       .mem_dqs_n
		memory_mem_odt     : out   std_logic;                                        --       .mem_odt
		memory_mem_dm      : out   std_logic_vector(3 downto 0);                     --       .mem_dm
		memory_oct_rzqin   : in    std_logic                     := '0';             --       .oct_rzqin
		reset_reset_n      : in    std_logic                     := '0'              --  reset.reset_n
	);
end entity soc;

architecture rtl of soc is
	component soc_hps_0 is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			mem_a                    : out   std_logic_vector(14 downto 0);                    -- mem_a
			mem_ba                   : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck                   : out   std_logic;                                        -- mem_ck
			mem_ck_n                 : out   std_logic;                                        -- mem_ck_n
			mem_cke                  : out   std_logic;                                        -- mem_cke
			mem_cs_n                 : out   std_logic;                                        -- mem_cs_n
			mem_ras_n                : out   std_logic;                                        -- mem_ras_n
			mem_cas_n                : out   std_logic;                                        -- mem_cas_n
			mem_we_n                 : out   std_logic;                                        -- mem_we_n
			mem_reset_n              : out   std_logic;                                        -- mem_reset_n
			mem_dq                   : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                  : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n                : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt                  : out   std_logic;                                        -- mem_odt
			mem_dm                   : out   std_logic_vector(3 downto 0);                     -- mem_dm
			oct_rzqin                : in    std_logic                     := 'X';             -- oct_rzqin
			h2f_rst_n                : out   std_logic;                                        -- reset_n
			f2h_sdram0_clk           : in    std_logic                     := 'X';             -- clk
			f2h_sdram0_ADDRESS       : in    std_logic_vector(28 downto 0) := (others => 'X'); -- address
			f2h_sdram0_BURSTCOUNT    : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- burstcount
			f2h_sdram0_WAITREQUEST   : out   std_logic;                                        -- waitrequest
			f2h_sdram0_WRITEDATA     : in    std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			f2h_sdram0_BYTEENABLE    : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			f2h_sdram0_WRITE         : in    std_logic                     := 'X';             -- write
			f2h_sdram1_clk           : in    std_logic                     := 'X';             -- clk
			f2h_sdram1_ADDRESS       : in    std_logic_vector(28 downto 0) := (others => 'X'); -- address
			f2h_sdram1_BURSTCOUNT    : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- burstcount
			f2h_sdram1_WAITREQUEST   : out   std_logic;                                        -- waitrequest
			f2h_sdram1_READDATA      : out   std_logic_vector(63 downto 0);                    -- readdata
			f2h_sdram1_READDATAVALID : out   std_logic;                                        -- readdatavalid
			f2h_sdram1_READ          : in    std_logic                     := 'X';             -- read
			h2f_lw_axi_clk           : in    std_logic                     := 'X';             -- clk
			h2f_lw_AWID              : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_lw_AWADDR            : out   std_logic_vector(20 downto 0);                    -- awaddr
			h2f_lw_AWLEN             : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_lw_AWSIZE            : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_lw_AWBURST           : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_lw_AWLOCK            : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_lw_AWCACHE           : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_lw_AWPROT            : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_lw_AWVALID           : out   std_logic;                                        -- awvalid
			h2f_lw_AWREADY           : in    std_logic                     := 'X';             -- awready
			h2f_lw_WID               : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_lw_WDATA             : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_lw_WSTRB             : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_lw_WLAST             : out   std_logic;                                        -- wlast
			h2f_lw_WVALID            : out   std_logic;                                        -- wvalid
			h2f_lw_WREADY            : in    std_logic                     := 'X';             -- wready
			h2f_lw_BID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_lw_BRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_lw_BVALID            : in    std_logic                     := 'X';             -- bvalid
			h2f_lw_BREADY            : out   std_logic;                                        -- bready
			h2f_lw_ARID              : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_lw_ARADDR            : out   std_logic_vector(20 downto 0);                    -- araddr
			h2f_lw_ARLEN             : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_lw_ARSIZE            : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_lw_ARBURST           : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_lw_ARLOCK            : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_lw_ARCACHE           : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_lw_ARPROT            : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_lw_ARVALID           : out   std_logic;                                        -- arvalid
			h2f_lw_ARREADY           : in    std_logic                     := 'X';             -- arready
			h2f_lw_RID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_lw_RDATA             : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_lw_RRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_lw_RLAST             : in    std_logic                     := 'X';             -- rlast
			h2f_lw_RVALID            : in    std_logic                     := 'X';             -- rvalid
			h2f_lw_RREADY            : out   std_logic                                         -- rready
		);
	end component soc_hps_0;

	component read_master is
		generic (
			DATA_WIDTH                : integer := 32;
			LENGTH_WIDTH              : integer := 32;
			FIFO_DEPTH                : integer := 32;
			STRIDE_ENABLE             : integer := 0;
			BURST_ENABLE              : integer := 0;
			PACKET_ENABLE             : integer := 0;
			ERROR_ENABLE              : integer := 0;
			ERROR_WIDTH               : integer := 8;
			CHANNEL_ENABLE            : integer := 0;
			CHANNEL_WIDTH             : integer := 8;
			BYTE_ENABLE_WIDTH         : integer := 4;
			BYTE_ENABLE_WIDTH_LOG2    : integer := 2;
			ADDRESS_WIDTH             : integer := 32;
			FIFO_DEPTH_LOG2           : integer := 5;
			SYMBOL_WIDTH              : integer := 8;
			NUMBER_OF_SYMBOLS         : integer := 4;
			NUMBER_OF_SYMBOLS_LOG2    : integer := 2;
			MAX_BURST_COUNT_WIDTH     : integer := 2;
			UNALIGNED_ACCESSES_ENABLE : integer := 0;
			ONLY_FULL_ACCESS_ENABLE   : integer := 0;
			BURST_WRAPPING_SUPPORT    : integer := 1;
			PROGRAMMABLE_BURST_ENABLE : integer := 0;
			MAX_BURST_COUNT           : integer := 2;
			FIFO_SPEED_OPTIMIZATION   : integer := 1;
			STRIDE_WIDTH              : integer := 1
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                     -- address
			master_read          : out std_logic;                                         -- read
			master_byteenable    : out std_logic_vector(7 downto 0);                      -- byteenable
			master_readdata      : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- readdata
			master_waitrequest   : in  std_logic                      := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                      := 'X';             -- readdatavalid
			src_data             : out std_logic_vector(63 downto 0);                     -- data
			src_valid            : out std_logic;                                         -- valid
			src_ready            : in  std_logic                      := 'X';             -- ready
			src_error            : out std_logic_vector(7 downto 0);                      -- error
			src_channel          : out std_logic_vector(7 downto 0);                      -- channel
			snk_command_data     : in  std_logic_vector(255 downto 0) := (others => 'X'); -- data
			snk_command_valid    : in  std_logic                      := 'X';             -- valid
			snk_command_ready    : out std_logic;                                         -- ready
			src_response_data    : out std_logic_vector(255 downto 0);                    -- data
			src_response_valid   : out std_logic;                                         -- valid
			src_response_ready   : in  std_logic                      := 'X';             -- ready
			master_burstcount    : out std_logic_vector(0 downto 0);                      -- burstcount
			src_sop              : out std_logic;                                         -- startofpacket
			src_eop              : out std_logic;                                         -- endofpacket
			src_empty            : out std_logic_vector(2 downto 0)                       -- empty
		);
	end component read_master;

	component altera_avalon_sc_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(63 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_error          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- error
			in_channel        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			out_data          : out std_logic_vector(63 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_error         : out std_logic_vector(7 downto 0);                     -- error
			out_channel       : out std_logic_vector(7 downto 0);                     -- channel
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic                                         -- empty
		);
	end component altera_avalon_sc_fifo;

	component write_master is
		generic (
			DATA_WIDTH                     : integer := 32;
			LENGTH_WIDTH                   : integer := 32;
			FIFO_DEPTH                     : integer := 32;
			STRIDE_ENABLE                  : integer := 0;
			BURST_ENABLE                   : integer := 0;
			PACKET_ENABLE                  : integer := 0;
			ERROR_ENABLE                   : integer := 0;
			ERROR_WIDTH                    : integer := 8;
			BYTE_ENABLE_WIDTH              : integer := 4;
			BYTE_ENABLE_WIDTH_LOG2         : integer := 2;
			ADDRESS_WIDTH                  : integer := 32;
			FIFO_DEPTH_LOG2                : integer := 5;
			SYMBOL_WIDTH                   : integer := 8;
			NUMBER_OF_SYMBOLS              : integer := 4;
			NUMBER_OF_SYMBOLS_LOG2         : integer := 2;
			MAX_BURST_COUNT_WIDTH          : integer := 2;
			UNALIGNED_ACCESSES_ENABLE      : integer := 0;
			ONLY_FULL_ACCESS_ENABLE        : integer := 0;
			BURST_WRAPPING_SUPPORT         : integer := 1;
			PROGRAMMABLE_BURST_ENABLE      : integer := 0;
			MAX_BURST_COUNT                : integer := 2;
			FIFO_SPEED_OPTIMIZATION        : integer := 1;
			STRIDE_WIDTH                   : integer := 1;
			ACTUAL_BYTES_TRANSFERRED_WIDTH : integer := 32
		);
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			master_address     : out std_logic_vector(31 downto 0);                     -- address
			master_write       : out std_logic;                                         -- write
			master_byteenable  : out std_logic_vector(7 downto 0);                      -- byteenable
			master_writedata   : out std_logic_vector(63 downto 0);                     -- writedata
			master_waitrequest : in  std_logic                      := 'X';             -- waitrequest
			snk_data           : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- data
			snk_valid          : in  std_logic                      := 'X';             -- valid
			snk_ready          : out std_logic;                                         -- ready
			snk_error          : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- error
			snk_command_data   : in  std_logic_vector(255 downto 0) := (others => 'X'); -- data
			snk_command_valid  : in  std_logic                      := 'X';             -- valid
			snk_command_ready  : out std_logic;                                         -- ready
			src_response_data  : out std_logic_vector(255 downto 0);                    -- data
			src_response_valid : out std_logic;                                         -- valid
			src_response_ready : in  std_logic                      := 'X';             -- ready
			master_burstcount  : out std_logic_vector(0 downto 0);                      -- burstcount
			snk_sop            : in  std_logic                      := 'X';             -- startofpacket
			snk_eop            : in  std_logic                      := 'X';             -- endofpacket
			snk_empty          : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- empty
		);
	end component write_master;

	component soc_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                                      : in  std_logic                     := 'X';             -- clk
			hps_0_f2h_sdram1_data_translator_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			read_master_sgdma_Clock_reset_reset_bridge_in_reset_reset          : in  std_logic                     := 'X';             -- reset
			read_master_sgdma_Data_Read_Master_address                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			read_master_sgdma_Data_Read_Master_waitrequest                     : out std_logic;                                        -- waitrequest
			read_master_sgdma_Data_Read_Master_byteenable                      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			read_master_sgdma_Data_Read_Master_read                            : in  std_logic                     := 'X';             -- read
			read_master_sgdma_Data_Read_Master_readdata                        : out std_logic_vector(63 downto 0);                    -- readdata
			read_master_sgdma_Data_Read_Master_readdatavalid                   : out std_logic;                                        -- readdatavalid
			hps_0_f2h_sdram1_data_address                                      : out std_logic_vector(28 downto 0);                    -- address
			hps_0_f2h_sdram1_data_read                                         : out std_logic;                                        -- read
			hps_0_f2h_sdram1_data_readdata                                     : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			hps_0_f2h_sdram1_data_burstcount                                   : out std_logic_vector(7 downto 0);                     -- burstcount
			hps_0_f2h_sdram1_data_readdatavalid                                : in  std_logic                     := 'X';             -- readdatavalid
			hps_0_f2h_sdram1_data_waitrequest                                  : in  std_logic                     := 'X'              -- waitrequest
		);
	end component soc_mm_interconnect_0;

	component soc_mm_interconnect_1 is
		port (
			clk_0_clk_clk                                                      : in  std_logic                     := 'X';             -- clk
			hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			write_master_sgdma_Clock_reset_reset_bridge_in_reset_reset         : in  std_logic                     := 'X';             -- reset
			write_master_sgdma_Data_Write_Master_address                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			write_master_sgdma_Data_Write_Master_waitrequest                   : out std_logic;                                        -- waitrequest
			write_master_sgdma_Data_Write_Master_byteenable                    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			write_master_sgdma_Data_Write_Master_write                         : in  std_logic                     := 'X';             -- write
			write_master_sgdma_Data_Write_Master_writedata                     : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			hps_0_f2h_sdram0_data_address                                      : out std_logic_vector(28 downto 0);                    -- address
			hps_0_f2h_sdram0_data_write                                        : out std_logic;                                        -- write
			hps_0_f2h_sdram0_data_writedata                                    : out std_logic_vector(63 downto 0);                    -- writedata
			hps_0_f2h_sdram0_data_burstcount                                   : out std_logic_vector(7 downto 0);                     -- burstcount
			hps_0_f2h_sdram0_data_byteenable                                   : out std_logic_vector(7 downto 0);                     -- byteenable
			hps_0_f2h_sdram0_data_waitrequest                                  : in  std_logic                     := 'X'              -- waitrequest
		);
	end component soc_mm_interconnect_1;

	component soc_mm_interconnect_2 is
		port (
			hps_0_h2f_lw_axi_master_awid                                        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- awid
			hps_0_h2f_lw_axi_master_awaddr                                      : in  std_logic_vector(20 downto 0)  := (others => 'X'); -- awaddr
			hps_0_h2f_lw_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awlen
			hps_0_h2f_lw_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awsize
			hps_0_h2f_lw_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- awburst
			hps_0_h2f_lw_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- awlock
			hps_0_h2f_lw_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awcache
			hps_0_h2f_lw_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awprot
			hps_0_h2f_lw_axi_master_awvalid                                     : in  std_logic                      := 'X';             -- awvalid
			hps_0_h2f_lw_axi_master_awready                                     : out std_logic;                                         -- awready
			hps_0_h2f_lw_axi_master_wid                                         : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- wid
			hps_0_h2f_lw_axi_master_wdata                                       : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- wdata
			hps_0_h2f_lw_axi_master_wstrb                                       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- wstrb
			hps_0_h2f_lw_axi_master_wlast                                       : in  std_logic                      := 'X';             -- wlast
			hps_0_h2f_lw_axi_master_wvalid                                      : in  std_logic                      := 'X';             -- wvalid
			hps_0_h2f_lw_axi_master_wready                                      : out std_logic;                                         -- wready
			hps_0_h2f_lw_axi_master_bid                                         : out std_logic_vector(11 downto 0);                     -- bid
			hps_0_h2f_lw_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                      -- bresp
			hps_0_h2f_lw_axi_master_bvalid                                      : out std_logic;                                         -- bvalid
			hps_0_h2f_lw_axi_master_bready                                      : in  std_logic                      := 'X';             -- bready
			hps_0_h2f_lw_axi_master_arid                                        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- arid
			hps_0_h2f_lw_axi_master_araddr                                      : in  std_logic_vector(20 downto 0)  := (others => 'X'); -- araddr
			hps_0_h2f_lw_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arlen
			hps_0_h2f_lw_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arsize
			hps_0_h2f_lw_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- arburst
			hps_0_h2f_lw_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- arlock
			hps_0_h2f_lw_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arcache
			hps_0_h2f_lw_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arprot
			hps_0_h2f_lw_axi_master_arvalid                                     : in  std_logic                      := 'X';             -- arvalid
			hps_0_h2f_lw_axi_master_arready                                     : out std_logic;                                         -- arready
			hps_0_h2f_lw_axi_master_rid                                         : out std_logic_vector(11 downto 0);                     -- rid
			hps_0_h2f_lw_axi_master_rdata                                       : out std_logic_vector(31 downto 0);                     -- rdata
			hps_0_h2f_lw_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                      -- rresp
			hps_0_h2f_lw_axi_master_rlast                                       : out std_logic;                                         -- rlast
			hps_0_h2f_lw_axi_master_rvalid                                      : out std_logic;                                         -- rvalid
			hps_0_h2f_lw_axi_master_rready                                      : in  std_logic                      := 'X';             -- rready
			clk_0_clk_clk                                                       : in  std_logic                      := 'X';             -- clk
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			sgdma_write_clock_reset_reset_bridge_in_reset_reset                 : in  std_logic                      := 'X';             -- reset
			sgdma_read_CSR_address                                              : out std_logic_vector(2 downto 0);                      -- address
			sgdma_read_CSR_write                                                : out std_logic;                                         -- write
			sgdma_read_CSR_read                                                 : out std_logic;                                         -- read
			sgdma_read_CSR_readdata                                             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			sgdma_read_CSR_writedata                                            : out std_logic_vector(31 downto 0);                     -- writedata
			sgdma_read_CSR_byteenable                                           : out std_logic_vector(3 downto 0);                      -- byteenable
			sgdma_read_Descriptor_Slave_write                                   : out std_logic;                                         -- write
			sgdma_read_Descriptor_Slave_writedata                               : out std_logic_vector(127 downto 0);                    -- writedata
			sgdma_read_Descriptor_Slave_byteenable                              : out std_logic_vector(15 downto 0);                     -- byteenable
			sgdma_read_Descriptor_Slave_waitrequest                             : in  std_logic                      := 'X';             -- waitrequest
			sgdma_write_CSR_address                                             : out std_logic_vector(2 downto 0);                      -- address
			sgdma_write_CSR_write                                               : out std_logic;                                         -- write
			sgdma_write_CSR_read                                                : out std_logic;                                         -- read
			sgdma_write_CSR_readdata                                            : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			sgdma_write_CSR_writedata                                           : out std_logic_vector(31 downto 0);                     -- writedata
			sgdma_write_CSR_byteenable                                          : out std_logic_vector(3 downto 0);                      -- byteenable
			sgdma_write_Descriptor_Slave_write                                  : out std_logic;                                         -- write
			sgdma_write_Descriptor_Slave_writedata                              : out std_logic_vector(127 downto 0);                    -- writedata
			sgdma_write_Descriptor_Slave_byteenable                             : out std_logic_vector(15 downto 0);                     -- byteenable
			sgdma_write_Descriptor_Slave_waitrequest                            : in  std_logic                      := 'X'              -- waitrequest
		);
	end component soc_mm_interconnect_2;

	component soc_avalon_st_adapter is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk   : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset : in  std_logic                     := 'X';             -- reset
			in_0_data      : in  std_logic_vector(63 downto 0) := (others => 'X'); -- data
			in_0_valid     : in  std_logic                     := 'X';             -- valid
			in_0_ready     : out std_logic;                                        -- ready
			in_0_error     : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- error
			in_0_channel   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			out_0_data     : out std_logic_vector(63 downto 0);                    -- data
			out_0_valid    : out std_logic;                                        -- valid
			out_0_ready    : in  std_logic                     := 'X';             -- ready
			out_0_error    : out std_logic_vector(7 downto 0)                      -- error
		);
	end component soc_avalon_st_adapter;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	component soc_sgdma_read is
		generic (
			MODE                        : integer := 0;
			RESPONSE_PORT               : integer := 0;
			DESCRIPTOR_FIFO_DEPTH       : integer := 128;
			ENHANCED_FEATURES           : integer := 1;
			DESCRIPTOR_WIDTH            : integer := 256;
			DESCRIPTOR_BYTEENABLE_WIDTH : integer := 32
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			csr_writedata           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write               : in  std_logic                      := 'X';             -- write
			csr_byteenable          : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata            : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                : in  std_logic                      := 'X';             -- read
			csr_address             : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_write        : in  std_logic                      := 'X';             -- write
			descriptor_waitrequest  : out std_logic;                                         -- waitrequest
			descriptor_writedata    : in  std_logic_vector(127 downto 0) := (others => 'X'); -- writedata
			descriptor_byteenable   : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- byteenable
			src_read_master_data    : out std_logic_vector(255 downto 0);                    -- data
			src_read_master_valid   : out std_logic;                                         -- valid
			src_read_master_ready   : in  std_logic                      := 'X';             -- ready
			snk_read_master_data    : in  std_logic_vector(255 downto 0) := (others => 'X'); -- data
			snk_read_master_valid   : in  std_logic                      := 'X';             -- valid
			snk_read_master_ready   : out std_logic;                                         -- ready
			csr_irq                 : out std_logic;                                         -- irq
			src_response_data       : out std_logic_vector(255 downto 0);                    -- data
			src_response_valid      : out std_logic;                                         -- valid
			src_response_ready      : in  std_logic                      := 'X';             -- ready
			mm_response_waitrequest : out std_logic;                                         -- waitrequest
			mm_response_byteenable  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			mm_response_address     : in  std_logic                      := 'X';             -- address
			mm_response_readdata    : out std_logic_vector(31 downto 0);                     -- readdata
			mm_response_read        : in  std_logic                      := 'X';             -- read
			src_write_master_data   : out std_logic_vector(255 downto 0);                    -- data
			src_write_master_valid  : out std_logic;                                         -- valid
			src_write_master_ready  : in  std_logic                      := 'X';             -- ready
			snk_write_master_data   : in  std_logic_vector(255 downto 0) := (others => 'X'); -- data
			snk_write_master_valid  : in  std_logic                      := 'X';             -- valid
			snk_write_master_ready  : out std_logic                                          -- ready
		);
	end component soc_sgdma_read;

	component soc_sgdma_write is
		generic (
			MODE                        : integer := 0;
			RESPONSE_PORT               : integer := 0;
			DESCRIPTOR_FIFO_DEPTH       : integer := 128;
			ENHANCED_FEATURES           : integer := 1;
			DESCRIPTOR_WIDTH            : integer := 256;
			DESCRIPTOR_BYTEENABLE_WIDTH : integer := 32
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			csr_writedata           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write               : in  std_logic                      := 'X';             -- write
			csr_byteenable          : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata            : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                : in  std_logic                      := 'X';             -- read
			csr_address             : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_write        : in  std_logic                      := 'X';             -- write
			descriptor_waitrequest  : out std_logic;                                         -- waitrequest
			descriptor_writedata    : in  std_logic_vector(127 downto 0) := (others => 'X'); -- writedata
			descriptor_byteenable   : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- byteenable
			src_write_master_data   : out std_logic_vector(255 downto 0);                    -- data
			src_write_master_valid  : out std_logic;                                         -- valid
			src_write_master_ready  : in  std_logic                      := 'X';             -- ready
			snk_write_master_data   : in  std_logic_vector(255 downto 0) := (others => 'X'); -- data
			snk_write_master_valid  : in  std_logic                      := 'X';             -- valid
			snk_write_master_ready  : out std_logic;                                         -- ready
			csr_irq                 : out std_logic;                                         -- irq
			src_response_data       : out std_logic_vector(255 downto 0);                    -- data
			src_response_valid      : out std_logic;                                         -- valid
			src_response_ready      : in  std_logic                      := 'X';             -- ready
			mm_response_waitrequest : out std_logic;                                         -- waitrequest
			mm_response_byteenable  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			mm_response_address     : in  std_logic                      := 'X';             -- address
			mm_response_readdata    : out std_logic_vector(31 downto 0);                     -- readdata
			mm_response_read        : in  std_logic                      := 'X';             -- read
			src_read_master_data    : out std_logic_vector(255 downto 0);                    -- data
			src_read_master_valid   : out std_logic;                                         -- valid
			src_read_master_ready   : in  std_logic                      := 'X';             -- ready
			snk_read_master_data    : in  std_logic_vector(255 downto 0) := (others => 'X'); -- data
			snk_read_master_valid   : in  std_logic                      := 'X';             -- valid
			snk_read_master_ready   : out std_logic                                          -- ready
		);
	end component soc_sgdma_write;

	signal read_master_sgdma_data_source_valid                        : std_logic;                      -- read_master_sgdma:src_valid -> sc_fifo_0:in_valid
	signal read_master_sgdma_data_source_data                         : std_logic_vector(63 downto 0);  -- read_master_sgdma:src_data -> sc_fifo_0:in_data
	signal read_master_sgdma_data_source_ready                        : std_logic;                      -- sc_fifo_0:in_ready -> read_master_sgdma:src_ready
	signal read_master_sgdma_data_source_channel                      : std_logic_vector(7 downto 0);   -- read_master_sgdma:src_channel -> sc_fifo_0:in_channel
	signal read_master_sgdma_data_source_error                        : std_logic_vector(7 downto 0);   -- read_master_sgdma:src_error -> sc_fifo_0:in_error
	signal sgdma_read_read_command_source_valid                       : std_logic;                      -- sgdma_read:src_read_master_valid -> read_master_sgdma:snk_command_valid
	signal sgdma_read_read_command_source_data                        : std_logic_vector(255 downto 0); -- sgdma_read:src_read_master_data -> read_master_sgdma:snk_command_data
	signal sgdma_read_read_command_source_ready                       : std_logic;                      -- read_master_sgdma:snk_command_ready -> sgdma_read:src_read_master_ready
	signal read_master_sgdma_response_source_valid                    : std_logic;                      -- read_master_sgdma:src_response_valid -> sgdma_read:snk_read_master_valid
	signal read_master_sgdma_response_source_data                     : std_logic_vector(255 downto 0); -- read_master_sgdma:src_response_data -> sgdma_read:snk_read_master_data
	signal read_master_sgdma_response_source_ready                    : std_logic;                      -- sgdma_read:snk_read_master_ready -> read_master_sgdma:src_response_ready
	signal write_master_sgdma_response_source_valid                   : std_logic;                      -- write_master_sgdma:src_response_valid -> sgdma_write:snk_write_master_valid
	signal write_master_sgdma_response_source_data                    : std_logic_vector(255 downto 0); -- write_master_sgdma:src_response_data -> sgdma_write:snk_write_master_data
	signal write_master_sgdma_response_source_ready                   : std_logic;                      -- sgdma_write:snk_write_master_ready -> write_master_sgdma:src_response_ready
	signal sgdma_write_write_command_source_valid                     : std_logic;                      -- sgdma_write:src_write_master_valid -> write_master_sgdma:snk_command_valid
	signal sgdma_write_write_command_source_data                      : std_logic_vector(255 downto 0); -- sgdma_write:src_write_master_data -> write_master_sgdma:snk_command_data
	signal sgdma_write_write_command_source_ready                     : std_logic;                      -- write_master_sgdma:snk_command_ready -> sgdma_write:src_write_master_ready
	signal read_master_sgdma_data_read_master_readdata                : std_logic_vector(63 downto 0);  -- mm_interconnect_0:read_master_sgdma_Data_Read_Master_readdata -> read_master_sgdma:master_readdata
	signal read_master_sgdma_data_read_master_waitrequest             : std_logic;                      -- mm_interconnect_0:read_master_sgdma_Data_Read_Master_waitrequest -> read_master_sgdma:master_waitrequest
	signal read_master_sgdma_data_read_master_address                 : std_logic_vector(31 downto 0);  -- read_master_sgdma:master_address -> mm_interconnect_0:read_master_sgdma_Data_Read_Master_address
	signal read_master_sgdma_data_read_master_read                    : std_logic;                      -- read_master_sgdma:master_read -> mm_interconnect_0:read_master_sgdma_Data_Read_Master_read
	signal read_master_sgdma_data_read_master_byteenable              : std_logic_vector(7 downto 0);   -- read_master_sgdma:master_byteenable -> mm_interconnect_0:read_master_sgdma_Data_Read_Master_byteenable
	signal read_master_sgdma_data_read_master_readdatavalid           : std_logic;                      -- mm_interconnect_0:read_master_sgdma_Data_Read_Master_readdatavalid -> read_master_sgdma:master_readdatavalid
	signal mm_interconnect_0_hps_0_f2h_sdram1_data_readdata           : std_logic_vector(63 downto 0);  -- hps_0:f2h_sdram1_READDATA -> mm_interconnect_0:hps_0_f2h_sdram1_data_readdata
	signal mm_interconnect_0_hps_0_f2h_sdram1_data_waitrequest        : std_logic;                      -- hps_0:f2h_sdram1_WAITREQUEST -> mm_interconnect_0:hps_0_f2h_sdram1_data_waitrequest
	signal mm_interconnect_0_hps_0_f2h_sdram1_data_address            : std_logic_vector(28 downto 0);  -- mm_interconnect_0:hps_0_f2h_sdram1_data_address -> hps_0:f2h_sdram1_ADDRESS
	signal mm_interconnect_0_hps_0_f2h_sdram1_data_read               : std_logic;                      -- mm_interconnect_0:hps_0_f2h_sdram1_data_read -> hps_0:f2h_sdram1_READ
	signal mm_interconnect_0_hps_0_f2h_sdram1_data_readdatavalid      : std_logic;                      -- hps_0:f2h_sdram1_READDATAVALID -> mm_interconnect_0:hps_0_f2h_sdram1_data_readdatavalid
	signal mm_interconnect_0_hps_0_f2h_sdram1_data_burstcount         : std_logic_vector(7 downto 0);   -- mm_interconnect_0:hps_0_f2h_sdram1_data_burstcount -> hps_0:f2h_sdram1_BURSTCOUNT
	signal write_master_sgdma_data_write_master_waitrequest           : std_logic;                      -- mm_interconnect_1:write_master_sgdma_Data_Write_Master_waitrequest -> write_master_sgdma:master_waitrequest
	signal write_master_sgdma_data_write_master_address               : std_logic_vector(31 downto 0);  -- write_master_sgdma:master_address -> mm_interconnect_1:write_master_sgdma_Data_Write_Master_address
	signal write_master_sgdma_data_write_master_byteenable            : std_logic_vector(7 downto 0);   -- write_master_sgdma:master_byteenable -> mm_interconnect_1:write_master_sgdma_Data_Write_Master_byteenable
	signal write_master_sgdma_data_write_master_write                 : std_logic;                      -- write_master_sgdma:master_write -> mm_interconnect_1:write_master_sgdma_Data_Write_Master_write
	signal write_master_sgdma_data_write_master_writedata             : std_logic_vector(63 downto 0);  -- write_master_sgdma:master_writedata -> mm_interconnect_1:write_master_sgdma_Data_Write_Master_writedata
	signal mm_interconnect_1_hps_0_f2h_sdram0_data_waitrequest        : std_logic;                      -- hps_0:f2h_sdram0_WAITREQUEST -> mm_interconnect_1:hps_0_f2h_sdram0_data_waitrequest
	signal mm_interconnect_1_hps_0_f2h_sdram0_data_address            : std_logic_vector(28 downto 0);  -- mm_interconnect_1:hps_0_f2h_sdram0_data_address -> hps_0:f2h_sdram0_ADDRESS
	signal mm_interconnect_1_hps_0_f2h_sdram0_data_byteenable         : std_logic_vector(7 downto 0);   -- mm_interconnect_1:hps_0_f2h_sdram0_data_byteenable -> hps_0:f2h_sdram0_BYTEENABLE
	signal mm_interconnect_1_hps_0_f2h_sdram0_data_write              : std_logic;                      -- mm_interconnect_1:hps_0_f2h_sdram0_data_write -> hps_0:f2h_sdram0_WRITE
	signal mm_interconnect_1_hps_0_f2h_sdram0_data_writedata          : std_logic_vector(63 downto 0);  -- mm_interconnect_1:hps_0_f2h_sdram0_data_writedata -> hps_0:f2h_sdram0_WRITEDATA
	signal mm_interconnect_1_hps_0_f2h_sdram0_data_burstcount         : std_logic_vector(7 downto 0);   -- mm_interconnect_1:hps_0_f2h_sdram0_data_burstcount -> hps_0:f2h_sdram0_BURSTCOUNT
	signal hps_0_h2f_lw_axi_master_awburst                            : std_logic_vector(1 downto 0);   -- hps_0:h2f_lw_AWBURST -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awburst
	signal hps_0_h2f_lw_axi_master_arlen                              : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_ARLEN -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arlen
	signal hps_0_h2f_lw_axi_master_wstrb                              : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_WSTRB -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wstrb
	signal hps_0_h2f_lw_axi_master_wready                             : std_logic;                      -- mm_interconnect_2:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	signal hps_0_h2f_lw_axi_master_rid                                : std_logic_vector(11 downto 0);  -- mm_interconnect_2:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	signal hps_0_h2f_lw_axi_master_rready                             : std_logic;                      -- hps_0:h2f_lw_RREADY -> mm_interconnect_2:hps_0_h2f_lw_axi_master_rready
	signal hps_0_h2f_lw_axi_master_awlen                              : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_AWLEN -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awlen
	signal hps_0_h2f_lw_axi_master_wid                                : std_logic_vector(11 downto 0);  -- hps_0:h2f_lw_WID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wid
	signal hps_0_h2f_lw_axi_master_arcache                            : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_ARCACHE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arcache
	signal hps_0_h2f_lw_axi_master_wvalid                             : std_logic;                      -- hps_0:h2f_lw_WVALID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wvalid
	signal hps_0_h2f_lw_axi_master_araddr                             : std_logic_vector(20 downto 0);  -- hps_0:h2f_lw_ARADDR -> mm_interconnect_2:hps_0_h2f_lw_axi_master_araddr
	signal hps_0_h2f_lw_axi_master_arprot                             : std_logic_vector(2 downto 0);   -- hps_0:h2f_lw_ARPROT -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arprot
	signal hps_0_h2f_lw_axi_master_awprot                             : std_logic_vector(2 downto 0);   -- hps_0:h2f_lw_AWPROT -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awprot
	signal hps_0_h2f_lw_axi_master_wdata                              : std_logic_vector(31 downto 0);  -- hps_0:h2f_lw_WDATA -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wdata
	signal hps_0_h2f_lw_axi_master_arvalid                            : std_logic;                      -- hps_0:h2f_lw_ARVALID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arvalid
	signal hps_0_h2f_lw_axi_master_awcache                            : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_AWCACHE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awcache
	signal hps_0_h2f_lw_axi_master_arid                               : std_logic_vector(11 downto 0);  -- hps_0:h2f_lw_ARID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arid
	signal hps_0_h2f_lw_axi_master_arlock                             : std_logic_vector(1 downto 0);   -- hps_0:h2f_lw_ARLOCK -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arlock
	signal hps_0_h2f_lw_axi_master_awlock                             : std_logic_vector(1 downto 0);   -- hps_0:h2f_lw_AWLOCK -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awlock
	signal hps_0_h2f_lw_axi_master_awaddr                             : std_logic_vector(20 downto 0);  -- hps_0:h2f_lw_AWADDR -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awaddr
	signal hps_0_h2f_lw_axi_master_bresp                              : std_logic_vector(1 downto 0);   -- mm_interconnect_2:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	signal hps_0_h2f_lw_axi_master_arready                            : std_logic;                      -- mm_interconnect_2:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	signal hps_0_h2f_lw_axi_master_rdata                              : std_logic_vector(31 downto 0);  -- mm_interconnect_2:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	signal hps_0_h2f_lw_axi_master_awready                            : std_logic;                      -- mm_interconnect_2:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	signal hps_0_h2f_lw_axi_master_arburst                            : std_logic_vector(1 downto 0);   -- hps_0:h2f_lw_ARBURST -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arburst
	signal hps_0_h2f_lw_axi_master_arsize                             : std_logic_vector(2 downto 0);   -- hps_0:h2f_lw_ARSIZE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arsize
	signal hps_0_h2f_lw_axi_master_bready                             : std_logic;                      -- hps_0:h2f_lw_BREADY -> mm_interconnect_2:hps_0_h2f_lw_axi_master_bready
	signal hps_0_h2f_lw_axi_master_rlast                              : std_logic;                      -- mm_interconnect_2:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	signal hps_0_h2f_lw_axi_master_wlast                              : std_logic;                      -- hps_0:h2f_lw_WLAST -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wlast
	signal hps_0_h2f_lw_axi_master_rresp                              : std_logic_vector(1 downto 0);   -- mm_interconnect_2:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	signal hps_0_h2f_lw_axi_master_awid                               : std_logic_vector(11 downto 0);  -- hps_0:h2f_lw_AWID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awid
	signal hps_0_h2f_lw_axi_master_bid                                : std_logic_vector(11 downto 0);  -- mm_interconnect_2:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	signal hps_0_h2f_lw_axi_master_bvalid                             : std_logic;                      -- mm_interconnect_2:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	signal hps_0_h2f_lw_axi_master_awsize                             : std_logic_vector(2 downto 0);   -- hps_0:h2f_lw_AWSIZE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awsize
	signal hps_0_h2f_lw_axi_master_awvalid                            : std_logic;                      -- hps_0:h2f_lw_AWVALID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awvalid
	signal hps_0_h2f_lw_axi_master_rvalid                             : std_logic;                      -- mm_interconnect_2:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	signal mm_interconnect_2_sgdma_write_csr_readdata                 : std_logic_vector(31 downto 0);  -- sgdma_write:csr_readdata -> mm_interconnect_2:sgdma_write_CSR_readdata
	signal mm_interconnect_2_sgdma_write_csr_address                  : std_logic_vector(2 downto 0);   -- mm_interconnect_2:sgdma_write_CSR_address -> sgdma_write:csr_address
	signal mm_interconnect_2_sgdma_write_csr_read                     : std_logic;                      -- mm_interconnect_2:sgdma_write_CSR_read -> sgdma_write:csr_read
	signal mm_interconnect_2_sgdma_write_csr_byteenable               : std_logic_vector(3 downto 0);   -- mm_interconnect_2:sgdma_write_CSR_byteenable -> sgdma_write:csr_byteenable
	signal mm_interconnect_2_sgdma_write_csr_write                    : std_logic;                      -- mm_interconnect_2:sgdma_write_CSR_write -> sgdma_write:csr_write
	signal mm_interconnect_2_sgdma_write_csr_writedata                : std_logic_vector(31 downto 0);  -- mm_interconnect_2:sgdma_write_CSR_writedata -> sgdma_write:csr_writedata
	signal mm_interconnect_2_sgdma_read_csr_readdata                  : std_logic_vector(31 downto 0);  -- sgdma_read:csr_readdata -> mm_interconnect_2:sgdma_read_CSR_readdata
	signal mm_interconnect_2_sgdma_read_csr_address                   : std_logic_vector(2 downto 0);   -- mm_interconnect_2:sgdma_read_CSR_address -> sgdma_read:csr_address
	signal mm_interconnect_2_sgdma_read_csr_read                      : std_logic;                      -- mm_interconnect_2:sgdma_read_CSR_read -> sgdma_read:csr_read
	signal mm_interconnect_2_sgdma_read_csr_byteenable                : std_logic_vector(3 downto 0);   -- mm_interconnect_2:sgdma_read_CSR_byteenable -> sgdma_read:csr_byteenable
	signal mm_interconnect_2_sgdma_read_csr_write                     : std_logic;                      -- mm_interconnect_2:sgdma_read_CSR_write -> sgdma_read:csr_write
	signal mm_interconnect_2_sgdma_read_csr_writedata                 : std_logic_vector(31 downto 0);  -- mm_interconnect_2:sgdma_read_CSR_writedata -> sgdma_read:csr_writedata
	signal mm_interconnect_2_sgdma_write_descriptor_slave_waitrequest : std_logic;                      -- sgdma_write:descriptor_waitrequest -> mm_interconnect_2:sgdma_write_Descriptor_Slave_waitrequest
	signal mm_interconnect_2_sgdma_write_descriptor_slave_byteenable  : std_logic_vector(15 downto 0);  -- mm_interconnect_2:sgdma_write_Descriptor_Slave_byteenable -> sgdma_write:descriptor_byteenable
	signal mm_interconnect_2_sgdma_write_descriptor_slave_write       : std_logic;                      -- mm_interconnect_2:sgdma_write_Descriptor_Slave_write -> sgdma_write:descriptor_write
	signal mm_interconnect_2_sgdma_write_descriptor_slave_writedata   : std_logic_vector(127 downto 0); -- mm_interconnect_2:sgdma_write_Descriptor_Slave_writedata -> sgdma_write:descriptor_writedata
	signal mm_interconnect_2_sgdma_read_descriptor_slave_waitrequest  : std_logic;                      -- sgdma_read:descriptor_waitrequest -> mm_interconnect_2:sgdma_read_Descriptor_Slave_waitrequest
	signal mm_interconnect_2_sgdma_read_descriptor_slave_byteenable   : std_logic_vector(15 downto 0);  -- mm_interconnect_2:sgdma_read_Descriptor_Slave_byteenable -> sgdma_read:descriptor_byteenable
	signal mm_interconnect_2_sgdma_read_descriptor_slave_write        : std_logic;                      -- mm_interconnect_2:sgdma_read_Descriptor_Slave_write -> sgdma_read:descriptor_write
	signal mm_interconnect_2_sgdma_read_descriptor_slave_writedata    : std_logic_vector(127 downto 0); -- mm_interconnect_2:sgdma_read_Descriptor_Slave_writedata -> sgdma_read:descriptor_writedata
	signal sc_fifo_0_out_valid                                        : std_logic;                      -- sc_fifo_0:out_valid -> avalon_st_adapter:in_0_valid
	signal sc_fifo_0_out_data                                         : std_logic_vector(63 downto 0);  -- sc_fifo_0:out_data -> avalon_st_adapter:in_0_data
	signal sc_fifo_0_out_ready                                        : std_logic;                      -- avalon_st_adapter:in_0_ready -> sc_fifo_0:out_ready
	signal sc_fifo_0_out_channel                                      : std_logic_vector(7 downto 0);   -- sc_fifo_0:out_channel -> avalon_st_adapter:in_0_channel
	signal sc_fifo_0_out_error                                        : std_logic_vector(7 downto 0);   -- sc_fifo_0:out_error -> avalon_st_adapter:in_0_error
	signal avalon_st_adapter_out_0_valid                              : std_logic;                      -- avalon_st_adapter:out_0_valid -> write_master_sgdma:snk_valid
	signal avalon_st_adapter_out_0_data                               : std_logic_vector(63 downto 0);  -- avalon_st_adapter:out_0_data -> write_master_sgdma:snk_data
	signal avalon_st_adapter_out_0_ready                              : std_logic;                      -- write_master_sgdma:snk_ready -> avalon_st_adapter:out_0_ready
	signal avalon_st_adapter_out_0_error                              : std_logic_vector(7 downto 0);   -- avalon_st_adapter:out_0_error -> write_master_sgdma:snk_error
	signal rst_controller_reset_out_reset                             : std_logic;                      -- rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, mm_interconnect_0:read_master_sgdma_Clock_reset_reset_bridge_in_reset_reset, mm_interconnect_1:write_master_sgdma_Clock_reset_reset_bridge_in_reset_reset, mm_interconnect_2:sgdma_write_clock_reset_reset_bridge_in_reset_reset, read_master_sgdma:reset, sc_fifo_0:reset, sgdma_read:reset, sgdma_write:reset, write_master_sgdma:reset]
	signal rst_controller_001_reset_out_reset                         : std_logic;                      -- rst_controller_001:reset_out -> [mm_interconnect_0:hps_0_f2h_sdram1_data_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_2:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]
	signal hps_0_h2f_reset_reset                                      : std_logic;                      -- hps_0:h2f_rst_n -> hps_0_h2f_reset_reset:in
	signal reset_reset_n_ports_inv                                    : std_logic;                      -- reset_reset_n:inv -> rst_controller:reset_in0
	signal hps_0_h2f_reset_reset_ports_inv                            : std_logic;                      -- hps_0_h2f_reset_reset:inv -> rst_controller_001:reset_in0

begin

	hps_0 : component soc_hps_0
		generic map (
			F2S_Width => 0,
			S2F_Width => 0
		)
		port map (
			mem_a                    => memory_mem_a,                                          --            memory.mem_a
			mem_ba                   => memory_mem_ba,                                         --                  .mem_ba
			mem_ck                   => memory_mem_ck,                                         --                  .mem_ck
			mem_ck_n                 => memory_mem_ck_n,                                       --                  .mem_ck_n
			mem_cke                  => memory_mem_cke,                                        --                  .mem_cke
			mem_cs_n                 => memory_mem_cs_n,                                       --                  .mem_cs_n
			mem_ras_n                => memory_mem_ras_n,                                      --                  .mem_ras_n
			mem_cas_n                => memory_mem_cas_n,                                      --                  .mem_cas_n
			mem_we_n                 => memory_mem_we_n,                                       --                  .mem_we_n
			mem_reset_n              => memory_mem_reset_n,                                    --                  .mem_reset_n
			mem_dq                   => memory_mem_dq,                                         --                  .mem_dq
			mem_dqs                  => memory_mem_dqs,                                        --                  .mem_dqs
			mem_dqs_n                => memory_mem_dqs_n,                                      --                  .mem_dqs_n
			mem_odt                  => memory_mem_odt,                                        --                  .mem_odt
			mem_dm                   => memory_mem_dm,                                         --                  .mem_dm
			oct_rzqin                => memory_oct_rzqin,                                      --                  .oct_rzqin
			h2f_rst_n                => hps_0_h2f_reset_reset,                                 --         h2f_reset.reset_n
			f2h_sdram0_clk           => clk_clk,                                               --  f2h_sdram0_clock.clk
			f2h_sdram0_ADDRESS       => mm_interconnect_1_hps_0_f2h_sdram0_data_address,       --   f2h_sdram0_data.address
			f2h_sdram0_BURSTCOUNT    => mm_interconnect_1_hps_0_f2h_sdram0_data_burstcount,    --                  .burstcount
			f2h_sdram0_WAITREQUEST   => mm_interconnect_1_hps_0_f2h_sdram0_data_waitrequest,   --                  .waitrequest
			f2h_sdram0_WRITEDATA     => mm_interconnect_1_hps_0_f2h_sdram0_data_writedata,     --                  .writedata
			f2h_sdram0_BYTEENABLE    => mm_interconnect_1_hps_0_f2h_sdram0_data_byteenable,    --                  .byteenable
			f2h_sdram0_WRITE         => mm_interconnect_1_hps_0_f2h_sdram0_data_write,         --                  .write
			f2h_sdram1_clk           => clk_clk,                                               --  f2h_sdram1_clock.clk
			f2h_sdram1_ADDRESS       => mm_interconnect_0_hps_0_f2h_sdram1_data_address,       --   f2h_sdram1_data.address
			f2h_sdram1_BURSTCOUNT    => mm_interconnect_0_hps_0_f2h_sdram1_data_burstcount,    --                  .burstcount
			f2h_sdram1_WAITREQUEST   => mm_interconnect_0_hps_0_f2h_sdram1_data_waitrequest,   --                  .waitrequest
			f2h_sdram1_READDATA      => mm_interconnect_0_hps_0_f2h_sdram1_data_readdata,      --                  .readdata
			f2h_sdram1_READDATAVALID => mm_interconnect_0_hps_0_f2h_sdram1_data_readdatavalid, --                  .readdatavalid
			f2h_sdram1_READ          => mm_interconnect_0_hps_0_f2h_sdram1_data_read,          --                  .read
			h2f_lw_axi_clk           => clk_clk,                                               --  h2f_lw_axi_clock.clk
			h2f_lw_AWID              => hps_0_h2f_lw_axi_master_awid,                          -- h2f_lw_axi_master.awid
			h2f_lw_AWADDR            => hps_0_h2f_lw_axi_master_awaddr,                        --                  .awaddr
			h2f_lw_AWLEN             => hps_0_h2f_lw_axi_master_awlen,                         --                  .awlen
			h2f_lw_AWSIZE            => hps_0_h2f_lw_axi_master_awsize,                        --                  .awsize
			h2f_lw_AWBURST           => hps_0_h2f_lw_axi_master_awburst,                       --                  .awburst
			h2f_lw_AWLOCK            => hps_0_h2f_lw_axi_master_awlock,                        --                  .awlock
			h2f_lw_AWCACHE           => hps_0_h2f_lw_axi_master_awcache,                       --                  .awcache
			h2f_lw_AWPROT            => hps_0_h2f_lw_axi_master_awprot,                        --                  .awprot
			h2f_lw_AWVALID           => hps_0_h2f_lw_axi_master_awvalid,                       --                  .awvalid
			h2f_lw_AWREADY           => hps_0_h2f_lw_axi_master_awready,                       --                  .awready
			h2f_lw_WID               => hps_0_h2f_lw_axi_master_wid,                           --                  .wid
			h2f_lw_WDATA             => hps_0_h2f_lw_axi_master_wdata,                         --                  .wdata
			h2f_lw_WSTRB             => hps_0_h2f_lw_axi_master_wstrb,                         --                  .wstrb
			h2f_lw_WLAST             => hps_0_h2f_lw_axi_master_wlast,                         --                  .wlast
			h2f_lw_WVALID            => hps_0_h2f_lw_axi_master_wvalid,                        --                  .wvalid
			h2f_lw_WREADY            => hps_0_h2f_lw_axi_master_wready,                        --                  .wready
			h2f_lw_BID               => hps_0_h2f_lw_axi_master_bid,                           --                  .bid
			h2f_lw_BRESP             => hps_0_h2f_lw_axi_master_bresp,                         --                  .bresp
			h2f_lw_BVALID            => hps_0_h2f_lw_axi_master_bvalid,                        --                  .bvalid
			h2f_lw_BREADY            => hps_0_h2f_lw_axi_master_bready,                        --                  .bready
			h2f_lw_ARID              => hps_0_h2f_lw_axi_master_arid,                          --                  .arid
			h2f_lw_ARADDR            => hps_0_h2f_lw_axi_master_araddr,                        --                  .araddr
			h2f_lw_ARLEN             => hps_0_h2f_lw_axi_master_arlen,                         --                  .arlen
			h2f_lw_ARSIZE            => hps_0_h2f_lw_axi_master_arsize,                        --                  .arsize
			h2f_lw_ARBURST           => hps_0_h2f_lw_axi_master_arburst,                       --                  .arburst
			h2f_lw_ARLOCK            => hps_0_h2f_lw_axi_master_arlock,                        --                  .arlock
			h2f_lw_ARCACHE           => hps_0_h2f_lw_axi_master_arcache,                       --                  .arcache
			h2f_lw_ARPROT            => hps_0_h2f_lw_axi_master_arprot,                        --                  .arprot
			h2f_lw_ARVALID           => hps_0_h2f_lw_axi_master_arvalid,                       --                  .arvalid
			h2f_lw_ARREADY           => hps_0_h2f_lw_axi_master_arready,                       --                  .arready
			h2f_lw_RID               => hps_0_h2f_lw_axi_master_rid,                           --                  .rid
			h2f_lw_RDATA             => hps_0_h2f_lw_axi_master_rdata,                         --                  .rdata
			h2f_lw_RRESP             => hps_0_h2f_lw_axi_master_rresp,                         --                  .rresp
			h2f_lw_RLAST             => hps_0_h2f_lw_axi_master_rlast,                         --                  .rlast
			h2f_lw_RVALID            => hps_0_h2f_lw_axi_master_rvalid,                        --                  .rvalid
			h2f_lw_RREADY            => hps_0_h2f_lw_axi_master_rready                         --                  .rready
		);

	read_master_sgdma : component read_master
		generic map (
			DATA_WIDTH                => 64,
			LENGTH_WIDTH              => 32,
			FIFO_DEPTH                => 128,
			STRIDE_ENABLE             => 0,
			BURST_ENABLE              => 0,
			PACKET_ENABLE             => 0,
			ERROR_ENABLE              => 1,
			ERROR_WIDTH               => 8,
			CHANNEL_ENABLE            => 1,
			CHANNEL_WIDTH             => 8,
			BYTE_ENABLE_WIDTH         => 8,
			BYTE_ENABLE_WIDTH_LOG2    => 3,
			ADDRESS_WIDTH             => 32,
			FIFO_DEPTH_LOG2           => 7,
			SYMBOL_WIDTH              => 8,
			NUMBER_OF_SYMBOLS         => 8,
			NUMBER_OF_SYMBOLS_LOG2    => 3,
			MAX_BURST_COUNT_WIDTH     => 1,
			UNALIGNED_ACCESSES_ENABLE => 0,
			ONLY_FULL_ACCESS_ENABLE   => 0,
			BURST_WRAPPING_SUPPORT    => 0,
			PROGRAMMABLE_BURST_ENABLE => 0,
			MAX_BURST_COUNT           => 1,
			FIFO_SPEED_OPTIMIZATION   => 1,
			STRIDE_WIDTH              => 1
		)
		port map (
			clk                  => clk_clk,                                          --            Clock.clk
			reset                => rst_controller_reset_out_reset,                   --      Clock_reset.reset
			master_address       => read_master_sgdma_data_read_master_address,       -- Data_Read_Master.address
			master_read          => read_master_sgdma_data_read_master_read,          --                 .read
			master_byteenable    => read_master_sgdma_data_read_master_byteenable,    --                 .byteenable
			master_readdata      => read_master_sgdma_data_read_master_readdata,      --                 .readdata
			master_waitrequest   => read_master_sgdma_data_read_master_waitrequest,   --                 .waitrequest
			master_readdatavalid => read_master_sgdma_data_read_master_readdatavalid, --                 .readdatavalid
			src_data             => read_master_sgdma_data_source_data,               --      Data_Source.data
			src_valid            => read_master_sgdma_data_source_valid,              --                 .valid
			src_ready            => read_master_sgdma_data_source_ready,              --                 .ready
			src_error            => read_master_sgdma_data_source_error,              --                 .error
			src_channel          => read_master_sgdma_data_source_channel,            --                 .channel
			snk_command_data     => sgdma_read_read_command_source_data,              --     Command_Sink.data
			snk_command_valid    => sgdma_read_read_command_source_valid,             --                 .valid
			snk_command_ready    => sgdma_read_read_command_source_ready,             --                 .ready
			src_response_data    => read_master_sgdma_response_source_data,           --  Response_Source.data
			src_response_valid   => read_master_sgdma_response_source_valid,          --                 .valid
			src_response_ready   => read_master_sgdma_response_source_ready,          --                 .ready
			master_burstcount    => open,                                             --      (terminated)
			src_sop              => open,                                             --      (terminated)
			src_eop              => open,                                             --      (terminated)
			src_empty            => open                                              --      (terminated)
		);

	sc_fifo_0 : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 8,
			BITS_PER_SYMBOL     => 8,
			FIFO_DEPTH          => 256,
			CHANNEL_WIDTH       => 8,
			ERROR_WIDTH         => 8,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 3,
			USE_MEMORY_BLOCKS   => 1,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                               --       clk.clk
			reset             => rst_controller_reset_out_reset,        -- clk_reset.reset
			in_data           => read_master_sgdma_data_source_data,    --        in.data
			in_valid          => read_master_sgdma_data_source_valid,   --          .valid
			in_ready          => read_master_sgdma_data_source_ready,   --          .ready
			in_error          => read_master_sgdma_data_source_error,   --          .error
			in_channel        => read_master_sgdma_data_source_channel, --          .channel
			out_data          => sc_fifo_0_out_data,                    --       out.data
			out_valid         => sc_fifo_0_out_valid,                   --          .valid
			out_ready         => sc_fifo_0_out_ready,                   --          .ready
			out_error         => sc_fifo_0_out_error,                   --          .error
			out_channel       => sc_fifo_0_out_channel,                 --          .channel
			csr_address       => "00",                                  -- (terminated)
			csr_read          => '0',                                   -- (terminated)
			csr_write         => '0',                                   -- (terminated)
			csr_readdata      => open,                                  -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",    -- (terminated)
			almost_full_data  => open,                                  -- (terminated)
			almost_empty_data => open,                                  -- (terminated)
			in_startofpacket  => '0',                                   -- (terminated)
			in_endofpacket    => '0',                                   -- (terminated)
			out_startofpacket => open,                                  -- (terminated)
			out_endofpacket   => open,                                  -- (terminated)
			in_empty          => '0',                                   -- (terminated)
			out_empty         => open                                   -- (terminated)
		);

	sgdma_read : component soc_sgdma_read
		generic map (
			MODE                        => 1,
			RESPONSE_PORT               => 2,
			DESCRIPTOR_FIFO_DEPTH       => 8,
			ENHANCED_FEATURES           => 0,
			DESCRIPTOR_WIDTH            => 128,
			DESCRIPTOR_BYTEENABLE_WIDTH => 16
		)
		port map (
			clk                     => clk_clk,                                                                                                                                                                                                                                                            --               clock.clk
			reset                   => rst_controller_reset_out_reset,                                                                                                                                                                                                                                     --         clock_reset.reset
			csr_writedata           => mm_interconnect_2_sgdma_read_csr_writedata,                                                                                                                                                                                                                         --                 CSR.writedata
			csr_write               => mm_interconnect_2_sgdma_read_csr_write,                                                                                                                                                                                                                             --                    .write
			csr_byteenable          => mm_interconnect_2_sgdma_read_csr_byteenable,                                                                                                                                                                                                                        --                    .byteenable
			csr_readdata            => mm_interconnect_2_sgdma_read_csr_readdata,                                                                                                                                                                                                                          --                    .readdata
			csr_read                => mm_interconnect_2_sgdma_read_csr_read,                                                                                                                                                                                                                              --                    .read
			csr_address             => mm_interconnect_2_sgdma_read_csr_address,                                                                                                                                                                                                                           --                    .address
			descriptor_write        => mm_interconnect_2_sgdma_read_descriptor_slave_write,                                                                                                                                                                                                                --    Descriptor_Slave.write
			descriptor_waitrequest  => mm_interconnect_2_sgdma_read_descriptor_slave_waitrequest,                                                                                                                                                                                                          --                    .waitrequest
			descriptor_writedata    => mm_interconnect_2_sgdma_read_descriptor_slave_writedata,                                                                                                                                                                                                            --                    .writedata
			descriptor_byteenable   => mm_interconnect_2_sgdma_read_descriptor_slave_byteenable,                                                                                                                                                                                                           --                    .byteenable
			src_read_master_data    => sgdma_read_read_command_source_data,                                                                                                                                                                                                                                -- Read_Command_Source.data
			src_read_master_valid   => sgdma_read_read_command_source_valid,                                                                                                                                                                                                                               --                    .valid
			src_read_master_ready   => sgdma_read_read_command_source_ready,                                                                                                                                                                                                                               --                    .ready
			snk_read_master_data    => read_master_sgdma_response_source_data,                                                                                                                                                                                                                             --  Read_Response_Sink.data
			snk_read_master_valid   => read_master_sgdma_response_source_valid,                                                                                                                                                                                                                            --                    .valid
			snk_read_master_ready   => read_master_sgdma_response_source_ready,                                                                                                                                                                                                                            --                    .ready
			csr_irq                 => open,                                                                                                                                                                                                                                                               --             csr_irq.irq
			src_response_data       => open,                                                                                                                                                                                                                                                               --         (terminated)
			src_response_valid      => open,                                                                                                                                                                                                                                                               --         (terminated)
			src_response_ready      => '0',                                                                                                                                                                                                                                                                --         (terminated)
			mm_response_waitrequest => open,                                                                                                                                                                                                                                                               --         (terminated)
			mm_response_byteenable  => "0000",                                                                                                                                                                                                                                                             --         (terminated)
			mm_response_address     => '0',                                                                                                                                                                                                                                                                --         (terminated)
			mm_response_readdata    => open,                                                                                                                                                                                                                                                               --         (terminated)
			mm_response_read        => '0',                                                                                                                                                                                                                                                                --         (terminated)
			src_write_master_data   => open,                                                                                                                                                                                                                                                               --         (terminated)
			src_write_master_valid  => open,                                                                                                                                                                                                                                                               --         (terminated)
			src_write_master_ready  => '0',                                                                                                                                                                                                                                                                --         (terminated)
			snk_write_master_data   => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --         (terminated)
			snk_write_master_valid  => '0',                                                                                                                                                                                                                                                                --         (terminated)
			snk_write_master_ready  => open                                                                                                                                                                                                                                                                --         (terminated)
		);

	sgdma_write : component soc_sgdma_write
		generic map (
			MODE                        => 2,
			RESPONSE_PORT               => 2,
			DESCRIPTOR_FIFO_DEPTH       => 8,
			ENHANCED_FEATURES           => 0,
			DESCRIPTOR_WIDTH            => 128,
			DESCRIPTOR_BYTEENABLE_WIDTH => 16
		)
		port map (
			clk                     => clk_clk,                                                                                                                                                                                                                                                            --                clock.clk
			reset                   => rst_controller_reset_out_reset,                                                                                                                                                                                                                                     --          clock_reset.reset
			csr_writedata           => mm_interconnect_2_sgdma_write_csr_writedata,                                                                                                                                                                                                                        --                  CSR.writedata
			csr_write               => mm_interconnect_2_sgdma_write_csr_write,                                                                                                                                                                                                                            --                     .write
			csr_byteenable          => mm_interconnect_2_sgdma_write_csr_byteenable,                                                                                                                                                                                                                       --                     .byteenable
			csr_readdata            => mm_interconnect_2_sgdma_write_csr_readdata,                                                                                                                                                                                                                         --                     .readdata
			csr_read                => mm_interconnect_2_sgdma_write_csr_read,                                                                                                                                                                                                                             --                     .read
			csr_address             => mm_interconnect_2_sgdma_write_csr_address,                                                                                                                                                                                                                          --                     .address
			descriptor_write        => mm_interconnect_2_sgdma_write_descriptor_slave_write,                                                                                                                                                                                                               --     Descriptor_Slave.write
			descriptor_waitrequest  => mm_interconnect_2_sgdma_write_descriptor_slave_waitrequest,                                                                                                                                                                                                         --                     .waitrequest
			descriptor_writedata    => mm_interconnect_2_sgdma_write_descriptor_slave_writedata,                                                                                                                                                                                                           --                     .writedata
			descriptor_byteenable   => mm_interconnect_2_sgdma_write_descriptor_slave_byteenable,                                                                                                                                                                                                          --                     .byteenable
			src_write_master_data   => sgdma_write_write_command_source_data,                                                                                                                                                                                                                              -- Write_Command_Source.data
			src_write_master_valid  => sgdma_write_write_command_source_valid,                                                                                                                                                                                                                             --                     .valid
			src_write_master_ready  => sgdma_write_write_command_source_ready,                                                                                                                                                                                                                             --                     .ready
			snk_write_master_data   => write_master_sgdma_response_source_data,                                                                                                                                                                                                                            --  Write_Response_Sink.data
			snk_write_master_valid  => write_master_sgdma_response_source_valid,                                                                                                                                                                                                                           --                     .valid
			snk_write_master_ready  => write_master_sgdma_response_source_ready,                                                                                                                                                                                                                           --                     .ready
			csr_irq                 => open,                                                                                                                                                                                                                                                               --              csr_irq.irq
			src_response_data       => open,                                                                                                                                                                                                                                                               --          (terminated)
			src_response_valid      => open,                                                                                                                                                                                                                                                               --          (terminated)
			src_response_ready      => '0',                                                                                                                                                                                                                                                                --          (terminated)
			mm_response_waitrequest => open,                                                                                                                                                                                                                                                               --          (terminated)
			mm_response_byteenable  => "0000",                                                                                                                                                                                                                                                             --          (terminated)
			mm_response_address     => '0',                                                                                                                                                                                                                                                                --          (terminated)
			mm_response_readdata    => open,                                                                                                                                                                                                                                                               --          (terminated)
			mm_response_read        => '0',                                                                                                                                                                                                                                                                --          (terminated)
			src_read_master_data    => open,                                                                                                                                                                                                                                                               --          (terminated)
			src_read_master_valid   => open,                                                                                                                                                                                                                                                               --          (terminated)
			src_read_master_ready   => '0',                                                                                                                                                                                                                                                                --          (terminated)
			snk_read_master_data    => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --          (terminated)
			snk_read_master_valid   => '0',                                                                                                                                                                                                                                                                --          (terminated)
			snk_read_master_ready   => open                                                                                                                                                                                                                                                                --          (terminated)
		);

	write_master_sgdma : component write_master
		generic map (
			DATA_WIDTH                     => 64,
			LENGTH_WIDTH                   => 32,
			FIFO_DEPTH                     => 128,
			STRIDE_ENABLE                  => 0,
			BURST_ENABLE                   => 0,
			PACKET_ENABLE                  => 0,
			ERROR_ENABLE                   => 1,
			ERROR_WIDTH                    => 8,
			BYTE_ENABLE_WIDTH              => 8,
			BYTE_ENABLE_WIDTH_LOG2         => 3,
			ADDRESS_WIDTH                  => 32,
			FIFO_DEPTH_LOG2                => 7,
			SYMBOL_WIDTH                   => 8,
			NUMBER_OF_SYMBOLS              => 8,
			NUMBER_OF_SYMBOLS_LOG2         => 3,
			MAX_BURST_COUNT_WIDTH          => 1,
			UNALIGNED_ACCESSES_ENABLE      => 0,
			ONLY_FULL_ACCESS_ENABLE        => 0,
			BURST_WRAPPING_SUPPORT         => 0,
			PROGRAMMABLE_BURST_ENABLE      => 0,
			MAX_BURST_COUNT                => 1,
			FIFO_SPEED_OPTIMIZATION        => 1,
			STRIDE_WIDTH                   => 1,
			ACTUAL_BYTES_TRANSFERRED_WIDTH => 32
		)
		port map (
			clk                => clk_clk,                                          --             Clock.clk
			reset              => rst_controller_reset_out_reset,                   --       Clock_reset.reset
			master_address     => write_master_sgdma_data_write_master_address,     -- Data_Write_Master.address
			master_write       => write_master_sgdma_data_write_master_write,       --                  .write
			master_byteenable  => write_master_sgdma_data_write_master_byteenable,  --                  .byteenable
			master_writedata   => write_master_sgdma_data_write_master_writedata,   --                  .writedata
			master_waitrequest => write_master_sgdma_data_write_master_waitrequest, --                  .waitrequest
			snk_data           => avalon_st_adapter_out_0_data,                     --         Data_Sink.data
			snk_valid          => avalon_st_adapter_out_0_valid,                    --                  .valid
			snk_ready          => avalon_st_adapter_out_0_ready,                    --                  .ready
			snk_error          => avalon_st_adapter_out_0_error,                    --                  .error
			snk_command_data   => sgdma_write_write_command_source_data,            --      Command_Sink.data
			snk_command_valid  => sgdma_write_write_command_source_valid,           --                  .valid
			snk_command_ready  => sgdma_write_write_command_source_ready,           --                  .ready
			src_response_data  => write_master_sgdma_response_source_data,          --   Response_Source.data
			src_response_valid => write_master_sgdma_response_source_valid,         --                  .valid
			src_response_ready => write_master_sgdma_response_source_ready,         --                  .ready
			master_burstcount  => open,                                             --       (terminated)
			snk_sop            => '0',                                              --       (terminated)
			snk_eop            => '0',                                              --       (terminated)
			snk_empty          => "000"                                             --       (terminated)
		);

	mm_interconnect_0 : component soc_mm_interconnect_0
		port map (
			clk_0_clk_clk                                                      => clk_clk,                                               --                                                    clk_0_clk.clk
			hps_0_f2h_sdram1_data_translator_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                    -- hps_0_f2h_sdram1_data_translator_reset_reset_bridge_in_reset.reset
			read_master_sgdma_Clock_reset_reset_bridge_in_reset_reset          => rst_controller_reset_out_reset,                        --          read_master_sgdma_Clock_reset_reset_bridge_in_reset.reset
			read_master_sgdma_Data_Read_Master_address                         => read_master_sgdma_data_read_master_address,            --                           read_master_sgdma_Data_Read_Master.address
			read_master_sgdma_Data_Read_Master_waitrequest                     => read_master_sgdma_data_read_master_waitrequest,        --                                                             .waitrequest
			read_master_sgdma_Data_Read_Master_byteenable                      => read_master_sgdma_data_read_master_byteenable,         --                                                             .byteenable
			read_master_sgdma_Data_Read_Master_read                            => read_master_sgdma_data_read_master_read,               --                                                             .read
			read_master_sgdma_Data_Read_Master_readdata                        => read_master_sgdma_data_read_master_readdata,           --                                                             .readdata
			read_master_sgdma_Data_Read_Master_readdatavalid                   => read_master_sgdma_data_read_master_readdatavalid,      --                                                             .readdatavalid
			hps_0_f2h_sdram1_data_address                                      => mm_interconnect_0_hps_0_f2h_sdram1_data_address,       --                                        hps_0_f2h_sdram1_data.address
			hps_0_f2h_sdram1_data_read                                         => mm_interconnect_0_hps_0_f2h_sdram1_data_read,          --                                                             .read
			hps_0_f2h_sdram1_data_readdata                                     => mm_interconnect_0_hps_0_f2h_sdram1_data_readdata,      --                                                             .readdata
			hps_0_f2h_sdram1_data_burstcount                                   => mm_interconnect_0_hps_0_f2h_sdram1_data_burstcount,    --                                                             .burstcount
			hps_0_f2h_sdram1_data_readdatavalid                                => mm_interconnect_0_hps_0_f2h_sdram1_data_readdatavalid, --                                                             .readdatavalid
			hps_0_f2h_sdram1_data_waitrequest                                  => mm_interconnect_0_hps_0_f2h_sdram1_data_waitrequest    --                                                             .waitrequest
		);

	mm_interconnect_1 : component soc_mm_interconnect_1
		port map (
			clk_0_clk_clk                                                      => clk_clk,                                             --                                                    clk_0_clk.clk
			hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                  -- hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset.reset
			write_master_sgdma_Clock_reset_reset_bridge_in_reset_reset         => rst_controller_reset_out_reset,                      --         write_master_sgdma_Clock_reset_reset_bridge_in_reset.reset
			write_master_sgdma_Data_Write_Master_address                       => write_master_sgdma_data_write_master_address,        --                         write_master_sgdma_Data_Write_Master.address
			write_master_sgdma_Data_Write_Master_waitrequest                   => write_master_sgdma_data_write_master_waitrequest,    --                                                             .waitrequest
			write_master_sgdma_Data_Write_Master_byteenable                    => write_master_sgdma_data_write_master_byteenable,     --                                                             .byteenable
			write_master_sgdma_Data_Write_Master_write                         => write_master_sgdma_data_write_master_write,          --                                                             .write
			write_master_sgdma_Data_Write_Master_writedata                     => write_master_sgdma_data_write_master_writedata,      --                                                             .writedata
			hps_0_f2h_sdram0_data_address                                      => mm_interconnect_1_hps_0_f2h_sdram0_data_address,     --                                        hps_0_f2h_sdram0_data.address
			hps_0_f2h_sdram0_data_write                                        => mm_interconnect_1_hps_0_f2h_sdram0_data_write,       --                                                             .write
			hps_0_f2h_sdram0_data_writedata                                    => mm_interconnect_1_hps_0_f2h_sdram0_data_writedata,   --                                                             .writedata
			hps_0_f2h_sdram0_data_burstcount                                   => mm_interconnect_1_hps_0_f2h_sdram0_data_burstcount,  --                                                             .burstcount
			hps_0_f2h_sdram0_data_byteenable                                   => mm_interconnect_1_hps_0_f2h_sdram0_data_byteenable,  --                                                             .byteenable
			hps_0_f2h_sdram0_data_waitrequest                                  => mm_interconnect_1_hps_0_f2h_sdram0_data_waitrequest  --                                                             .waitrequest
		);

	mm_interconnect_2 : component soc_mm_interconnect_2
		port map (
			hps_0_h2f_lw_axi_master_awid                                        => hps_0_h2f_lw_axi_master_awid,                               --                                       hps_0_h2f_lw_axi_master.awid
			hps_0_h2f_lw_axi_master_awaddr                                      => hps_0_h2f_lw_axi_master_awaddr,                             --                                                              .awaddr
			hps_0_h2f_lw_axi_master_awlen                                       => hps_0_h2f_lw_axi_master_awlen,                              --                                                              .awlen
			hps_0_h2f_lw_axi_master_awsize                                      => hps_0_h2f_lw_axi_master_awsize,                             --                                                              .awsize
			hps_0_h2f_lw_axi_master_awburst                                     => hps_0_h2f_lw_axi_master_awburst,                            --                                                              .awburst
			hps_0_h2f_lw_axi_master_awlock                                      => hps_0_h2f_lw_axi_master_awlock,                             --                                                              .awlock
			hps_0_h2f_lw_axi_master_awcache                                     => hps_0_h2f_lw_axi_master_awcache,                            --                                                              .awcache
			hps_0_h2f_lw_axi_master_awprot                                      => hps_0_h2f_lw_axi_master_awprot,                             --                                                              .awprot
			hps_0_h2f_lw_axi_master_awvalid                                     => hps_0_h2f_lw_axi_master_awvalid,                            --                                                              .awvalid
			hps_0_h2f_lw_axi_master_awready                                     => hps_0_h2f_lw_axi_master_awready,                            --                                                              .awready
			hps_0_h2f_lw_axi_master_wid                                         => hps_0_h2f_lw_axi_master_wid,                                --                                                              .wid
			hps_0_h2f_lw_axi_master_wdata                                       => hps_0_h2f_lw_axi_master_wdata,                              --                                                              .wdata
			hps_0_h2f_lw_axi_master_wstrb                                       => hps_0_h2f_lw_axi_master_wstrb,                              --                                                              .wstrb
			hps_0_h2f_lw_axi_master_wlast                                       => hps_0_h2f_lw_axi_master_wlast,                              --                                                              .wlast
			hps_0_h2f_lw_axi_master_wvalid                                      => hps_0_h2f_lw_axi_master_wvalid,                             --                                                              .wvalid
			hps_0_h2f_lw_axi_master_wready                                      => hps_0_h2f_lw_axi_master_wready,                             --                                                              .wready
			hps_0_h2f_lw_axi_master_bid                                         => hps_0_h2f_lw_axi_master_bid,                                --                                                              .bid
			hps_0_h2f_lw_axi_master_bresp                                       => hps_0_h2f_lw_axi_master_bresp,                              --                                                              .bresp
			hps_0_h2f_lw_axi_master_bvalid                                      => hps_0_h2f_lw_axi_master_bvalid,                             --                                                              .bvalid
			hps_0_h2f_lw_axi_master_bready                                      => hps_0_h2f_lw_axi_master_bready,                             --                                                              .bready
			hps_0_h2f_lw_axi_master_arid                                        => hps_0_h2f_lw_axi_master_arid,                               --                                                              .arid
			hps_0_h2f_lw_axi_master_araddr                                      => hps_0_h2f_lw_axi_master_araddr,                             --                                                              .araddr
			hps_0_h2f_lw_axi_master_arlen                                       => hps_0_h2f_lw_axi_master_arlen,                              --                                                              .arlen
			hps_0_h2f_lw_axi_master_arsize                                      => hps_0_h2f_lw_axi_master_arsize,                             --                                                              .arsize
			hps_0_h2f_lw_axi_master_arburst                                     => hps_0_h2f_lw_axi_master_arburst,                            --                                                              .arburst
			hps_0_h2f_lw_axi_master_arlock                                      => hps_0_h2f_lw_axi_master_arlock,                             --                                                              .arlock
			hps_0_h2f_lw_axi_master_arcache                                     => hps_0_h2f_lw_axi_master_arcache,                            --                                                              .arcache
			hps_0_h2f_lw_axi_master_arprot                                      => hps_0_h2f_lw_axi_master_arprot,                             --                                                              .arprot
			hps_0_h2f_lw_axi_master_arvalid                                     => hps_0_h2f_lw_axi_master_arvalid,                            --                                                              .arvalid
			hps_0_h2f_lw_axi_master_arready                                     => hps_0_h2f_lw_axi_master_arready,                            --                                                              .arready
			hps_0_h2f_lw_axi_master_rid                                         => hps_0_h2f_lw_axi_master_rid,                                --                                                              .rid
			hps_0_h2f_lw_axi_master_rdata                                       => hps_0_h2f_lw_axi_master_rdata,                              --                                                              .rdata
			hps_0_h2f_lw_axi_master_rresp                                       => hps_0_h2f_lw_axi_master_rresp,                              --                                                              .rresp
			hps_0_h2f_lw_axi_master_rlast                                       => hps_0_h2f_lw_axi_master_rlast,                              --                                                              .rlast
			hps_0_h2f_lw_axi_master_rvalid                                      => hps_0_h2f_lw_axi_master_rvalid,                             --                                                              .rvalid
			hps_0_h2f_lw_axi_master_rready                                      => hps_0_h2f_lw_axi_master_rready,                             --                                                              .rready
			clk_0_clk_clk                                                       => clk_clk,                                                    --                                                     clk_0_clk.clk
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                         -- hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			sgdma_write_clock_reset_reset_bridge_in_reset_reset                 => rst_controller_reset_out_reset,                             --                 sgdma_write_clock_reset_reset_bridge_in_reset.reset
			sgdma_read_CSR_address                                              => mm_interconnect_2_sgdma_read_csr_address,                   --                                                sgdma_read_CSR.address
			sgdma_read_CSR_write                                                => mm_interconnect_2_sgdma_read_csr_write,                     --                                                              .write
			sgdma_read_CSR_read                                                 => mm_interconnect_2_sgdma_read_csr_read,                      --                                                              .read
			sgdma_read_CSR_readdata                                             => mm_interconnect_2_sgdma_read_csr_readdata,                  --                                                              .readdata
			sgdma_read_CSR_writedata                                            => mm_interconnect_2_sgdma_read_csr_writedata,                 --                                                              .writedata
			sgdma_read_CSR_byteenable                                           => mm_interconnect_2_sgdma_read_csr_byteenable,                --                                                              .byteenable
			sgdma_read_Descriptor_Slave_write                                   => mm_interconnect_2_sgdma_read_descriptor_slave_write,        --                                   sgdma_read_Descriptor_Slave.write
			sgdma_read_Descriptor_Slave_writedata                               => mm_interconnect_2_sgdma_read_descriptor_slave_writedata,    --                                                              .writedata
			sgdma_read_Descriptor_Slave_byteenable                              => mm_interconnect_2_sgdma_read_descriptor_slave_byteenable,   --                                                              .byteenable
			sgdma_read_Descriptor_Slave_waitrequest                             => mm_interconnect_2_sgdma_read_descriptor_slave_waitrequest,  --                                                              .waitrequest
			sgdma_write_CSR_address                                             => mm_interconnect_2_sgdma_write_csr_address,                  --                                               sgdma_write_CSR.address
			sgdma_write_CSR_write                                               => mm_interconnect_2_sgdma_write_csr_write,                    --                                                              .write
			sgdma_write_CSR_read                                                => mm_interconnect_2_sgdma_write_csr_read,                     --                                                              .read
			sgdma_write_CSR_readdata                                            => mm_interconnect_2_sgdma_write_csr_readdata,                 --                                                              .readdata
			sgdma_write_CSR_writedata                                           => mm_interconnect_2_sgdma_write_csr_writedata,                --                                                              .writedata
			sgdma_write_CSR_byteenable                                          => mm_interconnect_2_sgdma_write_csr_byteenable,               --                                                              .byteenable
			sgdma_write_Descriptor_Slave_write                                  => mm_interconnect_2_sgdma_write_descriptor_slave_write,       --                                  sgdma_write_Descriptor_Slave.write
			sgdma_write_Descriptor_Slave_writedata                              => mm_interconnect_2_sgdma_write_descriptor_slave_writedata,   --                                                              .writedata
			sgdma_write_Descriptor_Slave_byteenable                             => mm_interconnect_2_sgdma_write_descriptor_slave_byteenable,  --                                                              .byteenable
			sgdma_write_Descriptor_Slave_waitrequest                            => mm_interconnect_2_sgdma_write_descriptor_slave_waitrequest  --                                                              .waitrequest
		);

	avalon_st_adapter : component soc_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 0,
			inDataWidth     => 64,
			inChannelWidth  => 8,
			inErrorWidth    => 8,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 64,
			outChannelWidth => 0,
			outErrorWidth   => 8,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk   => clk_clk,                        -- in_clk_0.clk
			in_rst_0_reset => rst_controller_reset_out_reset, -- in_rst_0.reset
			in_0_data      => sc_fifo_0_out_data,             --     in_0.data
			in_0_valid     => sc_fifo_0_out_valid,            --         .valid
			in_0_ready     => sc_fifo_0_out_ready,            --         .ready
			in_0_error     => sc_fifo_0_out_error,            --         .error
			in_0_channel   => sc_fifo_0_out_channel,          --         .channel
			out_0_data     => avalon_st_adapter_out_0_data,   --    out_0.data
			out_0_valid    => avalon_st_adapter_out_0_valid,  --         .valid
			out_0_ready    => avalon_st_adapter_out_0_ready,  --         .ready
			out_0_error    => avalon_st_adapter_out_0_error   --         .error
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_0_h2f_reset_reset_ports_inv,    -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	hps_0_h2f_reset_reset_ports_inv <= not hps_0_h2f_reset_reset;

end architecture rtl; -- of soc
