-- soc.vhd

-- Generated using ACDS version 15.0 145

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc is
	port (
		clk_clk            : in    std_logic                     := '0';             --        clk.clk
		memory_mem_a       : out   std_logic_vector(14 downto 0);                    --     memory.mem_a
		memory_mem_ba      : out   std_logic_vector(2 downto 0);                     --           .mem_ba
		memory_mem_ck      : out   std_logic;                                        --           .mem_ck
		memory_mem_ck_n    : out   std_logic;                                        --           .mem_ck_n
		memory_mem_cke     : out   std_logic;                                        --           .mem_cke
		memory_mem_cs_n    : out   std_logic;                                        --           .mem_cs_n
		memory_mem_ras_n   : out   std_logic;                                        --           .mem_ras_n
		memory_mem_cas_n   : out   std_logic;                                        --           .mem_cas_n
		memory_mem_we_n    : out   std_logic;                                        --           .mem_we_n
		memory_mem_reset_n : out   std_logic;                                        --           .mem_reset_n
		memory_mem_dq      : inout std_logic_vector(31 downto 0) := (others => '0'); --           .mem_dq
		memory_mem_dqs     : inout std_logic_vector(3 downto 0)  := (others => '0'); --           .mem_dqs
		memory_mem_dqs_n   : inout std_logic_vector(3 downto 0)  := (others => '0'); --           .mem_dqs_n
		memory_mem_odt     : out   std_logic;                                        --           .mem_odt
		memory_mem_dm      : out   std_logic_vector(3 downto 0);                     --           .mem_dm
		memory_oct_rzqin   : in    std_logic                     := '0';             --           .oct_rzqin
		reccontrol_enrec   : out   std_logic;                                        -- reccontrol.enrec
		reset_reset_n      : in    std_logic                     := '0';             --      reset.reset_n
		rfrec_rxclock      : in    std_logic                     := '0';             --      rfrec.rxclock
		rfrec_rxdata       : in    std_logic_vector(11 downto 0) := (others => '0'); --           .rxdata
		rfrec_rxenable     : out   std_logic;                                        --           .rxenable
		rfrec_rxiq         : in    std_logic                     := '0';             --           .rxiq
		rfrec_recen        : in    std_logic                     := '0';             --           .recen
		rfrec_testled      : out   std_logic_vector(3 downto 0)                      --           .testled
	);
end entity soc;

architecture rtl of soc is
	component altera_avalon_dc_fifo is
		generic (
			SYMBOLS_PER_BEAT   : integer := 1;
			BITS_PER_SYMBOL    : integer := 8;
			FIFO_DEPTH         : integer := 16;
			CHANNEL_WIDTH      : integer := 0;
			ERROR_WIDTH        : integer := 0;
			USE_PACKETS        : integer := 0;
			USE_IN_FILL_LEVEL  : integer := 0;
			USE_OUT_FILL_LEVEL : integer := 0;
			WR_SYNC_DEPTH      : integer := 3;
			RD_SYNC_DEPTH      : integer := 3
		);
		port (
			in_clk            : in  std_logic                     := 'X';             -- clk
			in_reset_n        : in  std_logic                     := 'X';             -- reset_n
			out_clk           : in  std_logic                     := 'X';             -- clk
			out_reset_n       : in  std_logic                     := 'X';             -- reset_n
			in_data           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			out_data          : out std_logic_vector(15 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			in_csr_address    : in  std_logic                     := 'X';             -- address
			in_csr_read       : in  std_logic                     := 'X';             -- read
			in_csr_write      : in  std_logic                     := 'X';             -- write
			in_csr_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_csr_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			out_csr_address   : in  std_logic                     := 'X';             -- address
			out_csr_read      : in  std_logic                     := 'X';             -- read
			out_csr_write     : in  std_logic                     := 'X';             -- write
			out_csr_readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			out_csr_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component altera_avalon_dc_fifo;

	component dispatcher is
		generic (
			MODE                        : integer := 0;
			RESPONSE_PORT               : integer := 0;
			DESCRIPTOR_FIFO_DEPTH       : integer := 128;
			ENHANCED_FEATURES           : integer := 1;
			DESCRIPTOR_WIDTH            : integer := 256;
			DESCRIPTOR_BYTEENABLE_WIDTH : integer := 32
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			csr_writedata           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write               : in  std_logic                      := 'X';             -- write
			csr_byteenable          : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata            : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                : in  std_logic                      := 'X';             -- read
			csr_address             : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_write        : in  std_logic                      := 'X';             -- write
			descriptor_waitrequest  : out std_logic;                                         -- waitrequest
			descriptor_writedata    : in  std_logic_vector(127 downto 0) := (others => 'X'); -- writedata
			descriptor_byteenable   : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- byteenable
			src_write_master_data   : out std_logic_vector(255 downto 0);                    -- data
			src_write_master_valid  : out std_logic;                                         -- valid
			src_write_master_ready  : in  std_logic                      := 'X';             -- ready
			snk_write_master_data   : in  std_logic_vector(255 downto 0) := (others => 'X'); -- data
			snk_write_master_valid  : in  std_logic                      := 'X';             -- valid
			snk_write_master_ready  : out std_logic;                                         -- ready
			csr_irq                 : out std_logic;                                         -- irq
			src_response_data       : out std_logic_vector(255 downto 0);                    -- data
			src_response_valid      : out std_logic;                                         -- valid
			src_response_ready      : in  std_logic                      := 'X';             -- ready
			mm_response_waitrequest : out std_logic;                                         -- waitrequest
			mm_response_byteenable  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			mm_response_address     : in  std_logic                      := 'X';             -- address
			mm_response_readdata    : out std_logic_vector(31 downto 0);                     -- readdata
			mm_response_read        : in  std_logic                      := 'X';             -- read
			src_read_master_data    : out std_logic_vector(255 downto 0);                    -- data
			src_read_master_valid   : out std_logic;                                         -- valid
			src_read_master_ready   : in  std_logic                      := 'X';             -- ready
			snk_read_master_data    : in  std_logic_vector(255 downto 0) := (others => 'X'); -- data
			snk_read_master_valid   : in  std_logic                      := 'X';             -- valid
			snk_read_master_ready   : out std_logic                                          -- ready
		);
	end component dispatcher;

	component write_master is
		generic (
			DATA_WIDTH                     : integer := 32;
			LENGTH_WIDTH                   : integer := 32;
			FIFO_DEPTH                     : integer := 32;
			STRIDE_ENABLE                  : integer := 0;
			BURST_ENABLE                   : integer := 0;
			PACKET_ENABLE                  : integer := 0;
			ERROR_ENABLE                   : integer := 0;
			ERROR_WIDTH                    : integer := 8;
			BYTE_ENABLE_WIDTH              : integer := 4;
			BYTE_ENABLE_WIDTH_LOG2         : integer := 2;
			ADDRESS_WIDTH                  : integer := 32;
			FIFO_DEPTH_LOG2                : integer := 5;
			SYMBOL_WIDTH                   : integer := 8;
			NUMBER_OF_SYMBOLS              : integer := 4;
			NUMBER_OF_SYMBOLS_LOG2         : integer := 2;
			MAX_BURST_COUNT_WIDTH          : integer := 2;
			UNALIGNED_ACCESSES_ENABLE      : integer := 0;
			ONLY_FULL_ACCESS_ENABLE        : integer := 0;
			BURST_WRAPPING_SUPPORT         : integer := 1;
			PROGRAMMABLE_BURST_ENABLE      : integer := 0;
			MAX_BURST_COUNT                : integer := 2;
			FIFO_SPEED_OPTIMIZATION        : integer := 1;
			STRIDE_WIDTH                   : integer := 1;
			ACTUAL_BYTES_TRANSFERRED_WIDTH : integer := 32
		);
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			master_address     : out std_logic_vector(31 downto 0);                     -- address
			master_write       : out std_logic;                                         -- write
			master_byteenable  : out std_logic_vector(1 downto 0);                      -- byteenable
			master_writedata   : out std_logic_vector(15 downto 0);                     -- writedata
			master_waitrequest : in  std_logic                      := 'X';             -- waitrequest
			snk_data           : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- data
			snk_valid          : in  std_logic                      := 'X';             -- valid
			snk_ready          : out std_logic;                                         -- ready
			snk_command_data   : in  std_logic_vector(255 downto 0) := (others => 'X'); -- data
			snk_command_valid  : in  std_logic                      := 'X';             -- valid
			snk_command_ready  : out std_logic;                                         -- ready
			src_response_data  : out std_logic_vector(255 downto 0);                    -- data
			src_response_valid : out std_logic;                                         -- valid
			src_response_ready : in  std_logic                      := 'X';             -- ready
			master_burstcount  : out std_logic_vector(0 downto 0);                      -- burstcount
			snk_sop            : in  std_logic                      := 'X';             -- startofpacket
			snk_eop            : in  std_logic                      := 'X';             -- endofpacket
			snk_empty          : in  std_logic                      := 'X';             -- empty
			snk_error          : in  std_logic_vector(7 downto 0)   := (others => 'X')  -- error
		);
	end component write_master;

	component RFReceive is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			RXCLK         : in  std_logic                     := 'X';             -- rxclock
			RXD           : in  std_logic_vector(11 downto 0) := (others => 'X'); -- rxdata
			RXEN          : out std_logic;                                        -- rxenable
			RXIQSEL       : in  std_logic                     := 'X';             -- rxiq
			RecEnable     : in  std_logic                     := 'X';             -- recen
			LED           : out std_logic_vector(3 downto 0);                     -- testled
			rfRec_i_data  : out std_logic_vector(15 downto 0);                    -- data
			rfRec_i_ready : in  std_logic                     := 'X';             -- ready
			rfRec_i_valid : out std_logic;                                        -- valid
			rfRec_q_data  : out std_logic_vector(15 downto 0);                    -- data
			rfRec_q_ready : in  std_logic                     := 'X';             -- ready
			rfRec_q_valid : out std_logic;                                        -- valid
			rfRec_i_clk   : out std_logic;                                        -- clk
			rfRec_q_clk   : out std_logic                                         -- clk
		);
	end component RFReceive;

	component soc_hps_0 is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			mem_a                  : out   std_logic_vector(14 downto 0);                    -- mem_a
			mem_ba                 : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck                 : out   std_logic;                                        -- mem_ck
			mem_ck_n               : out   std_logic;                                        -- mem_ck_n
			mem_cke                : out   std_logic;                                        -- mem_cke
			mem_cs_n               : out   std_logic;                                        -- mem_cs_n
			mem_ras_n              : out   std_logic;                                        -- mem_ras_n
			mem_cas_n              : out   std_logic;                                        -- mem_cas_n
			mem_we_n               : out   std_logic;                                        -- mem_we_n
			mem_reset_n            : out   std_logic;                                        -- mem_reset_n
			mem_dq                 : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n              : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt                : out   std_logic;                                        -- mem_odt
			mem_dm                 : out   std_logic_vector(3 downto 0);                     -- mem_dm
			oct_rzqin              : in    std_logic                     := 'X';             -- oct_rzqin
			h2f_rst_n              : out   std_logic;                                        -- reset_n
			f2h_sdram0_clk         : in    std_logic                     := 'X';             -- clk
			f2h_sdram0_ADDRESS     : in    std_logic_vector(28 downto 0) := (others => 'X'); -- address
			f2h_sdram0_BURSTCOUNT  : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- burstcount
			f2h_sdram0_WAITREQUEST : out   std_logic;                                        -- waitrequest
			f2h_sdram0_WRITEDATA   : in    std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			f2h_sdram0_BYTEENABLE  : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			f2h_sdram0_WRITE       : in    std_logic                     := 'X';             -- write
			h2f_lw_axi_clk         : in    std_logic                     := 'X';             -- clk
			h2f_lw_AWID            : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_lw_AWADDR          : out   std_logic_vector(20 downto 0);                    -- awaddr
			h2f_lw_AWLEN           : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_lw_AWSIZE          : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_lw_AWBURST         : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_lw_AWLOCK          : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_lw_AWCACHE         : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_lw_AWPROT          : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_lw_AWVALID         : out   std_logic;                                        -- awvalid
			h2f_lw_AWREADY         : in    std_logic                     := 'X';             -- awready
			h2f_lw_WID             : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_lw_WDATA           : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_lw_WSTRB           : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_lw_WLAST           : out   std_logic;                                        -- wlast
			h2f_lw_WVALID          : out   std_logic;                                        -- wvalid
			h2f_lw_WREADY          : in    std_logic                     := 'X';             -- wready
			h2f_lw_BID             : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_lw_BRESP           : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_lw_BVALID          : in    std_logic                     := 'X';             -- bvalid
			h2f_lw_BREADY          : out   std_logic;                                        -- bready
			h2f_lw_ARID            : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_lw_ARADDR          : out   std_logic_vector(20 downto 0);                    -- araddr
			h2f_lw_ARLEN           : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_lw_ARSIZE          : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_lw_ARBURST         : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_lw_ARLOCK          : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_lw_ARCACHE         : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_lw_ARPROT          : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_lw_ARVALID         : out   std_logic;                                        -- arvalid
			h2f_lw_ARREADY         : in    std_logic                     := 'X';             -- arready
			h2f_lw_RID             : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_lw_RDATA           : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_lw_RRESP           : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_lw_RLAST           : in    std_logic                     := 'X';             -- rlast
			h2f_lw_RVALID          : in    std_logic                     := 'X';             -- rvalid
			h2f_lw_RREADY          : out   std_logic                                         -- rready
		);
	end component soc_hps_0;

	component recCtrl is
		port (
			clk        : in  std_logic                    := 'X';             -- clk
			reset      : in  std_logic                    := 'X';             -- reset
			RecEnable  : out std_logic;                                       -- enrec
			write_data : in  std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			write_en   : in  std_logic                    := 'X'              -- write
		);
	end component recCtrl;

	component soc_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                                      : in  std_logic                     := 'X';             -- clk
			hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			IN_WRITE_MASTER_Clock_reset_reset_bridge_in_reset_reset            : in  std_logic                     := 'X';             -- reset
			IN_WRITE_MASTER_Data_Write_Master_address                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			IN_WRITE_MASTER_Data_Write_Master_waitrequest                      : out std_logic;                                        -- waitrequest
			IN_WRITE_MASTER_Data_Write_Master_byteenable                       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			IN_WRITE_MASTER_Data_Write_Master_write                            : in  std_logic                     := 'X';             -- write
			IN_WRITE_MASTER_Data_Write_Master_writedata                        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			QU_WRITE_MASTER_Data_Write_Master_address                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			QU_WRITE_MASTER_Data_Write_Master_waitrequest                      : out std_logic;                                        -- waitrequest
			QU_WRITE_MASTER_Data_Write_Master_byteenable                       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			QU_WRITE_MASTER_Data_Write_Master_write                            : in  std_logic                     := 'X';             -- write
			QU_WRITE_MASTER_Data_Write_Master_writedata                        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			hps_0_f2h_sdram0_data_address                                      : out std_logic_vector(28 downto 0);                    -- address
			hps_0_f2h_sdram0_data_write                                        : out std_logic;                                        -- write
			hps_0_f2h_sdram0_data_writedata                                    : out std_logic_vector(63 downto 0);                    -- writedata
			hps_0_f2h_sdram0_data_burstcount                                   : out std_logic_vector(7 downto 0);                     -- burstcount
			hps_0_f2h_sdram0_data_byteenable                                   : out std_logic_vector(7 downto 0);                     -- byteenable
			hps_0_f2h_sdram0_data_waitrequest                                  : in  std_logic                     := 'X'              -- waitrequest
		);
	end component soc_mm_interconnect_0;

	component soc_mm_interconnect_1 is
		port (
			hps_0_h2f_lw_axi_master_awid                                        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- awid
			hps_0_h2f_lw_axi_master_awaddr                                      : in  std_logic_vector(20 downto 0)  := (others => 'X'); -- awaddr
			hps_0_h2f_lw_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awlen
			hps_0_h2f_lw_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awsize
			hps_0_h2f_lw_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- awburst
			hps_0_h2f_lw_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- awlock
			hps_0_h2f_lw_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awcache
			hps_0_h2f_lw_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awprot
			hps_0_h2f_lw_axi_master_awvalid                                     : in  std_logic                      := 'X';             -- awvalid
			hps_0_h2f_lw_axi_master_awready                                     : out std_logic;                                         -- awready
			hps_0_h2f_lw_axi_master_wid                                         : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- wid
			hps_0_h2f_lw_axi_master_wdata                                       : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- wdata
			hps_0_h2f_lw_axi_master_wstrb                                       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- wstrb
			hps_0_h2f_lw_axi_master_wlast                                       : in  std_logic                      := 'X';             -- wlast
			hps_0_h2f_lw_axi_master_wvalid                                      : in  std_logic                      := 'X';             -- wvalid
			hps_0_h2f_lw_axi_master_wready                                      : out std_logic;                                         -- wready
			hps_0_h2f_lw_axi_master_bid                                         : out std_logic_vector(11 downto 0);                     -- bid
			hps_0_h2f_lw_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                      -- bresp
			hps_0_h2f_lw_axi_master_bvalid                                      : out std_logic;                                         -- bvalid
			hps_0_h2f_lw_axi_master_bready                                      : in  std_logic                      := 'X';             -- bready
			hps_0_h2f_lw_axi_master_arid                                        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- arid
			hps_0_h2f_lw_axi_master_araddr                                      : in  std_logic_vector(20 downto 0)  := (others => 'X'); -- araddr
			hps_0_h2f_lw_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arlen
			hps_0_h2f_lw_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arsize
			hps_0_h2f_lw_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- arburst
			hps_0_h2f_lw_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- arlock
			hps_0_h2f_lw_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arcache
			hps_0_h2f_lw_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arprot
			hps_0_h2f_lw_axi_master_arvalid                                     : in  std_logic                      := 'X';             -- arvalid
			hps_0_h2f_lw_axi_master_arready                                     : out std_logic;                                         -- arready
			hps_0_h2f_lw_axi_master_rid                                         : out std_logic_vector(11 downto 0);                     -- rid
			hps_0_h2f_lw_axi_master_rdata                                       : out std_logic_vector(31 downto 0);                     -- rdata
			hps_0_h2f_lw_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                      -- rresp
			hps_0_h2f_lw_axi_master_rlast                                       : out std_logic;                                         -- rlast
			hps_0_h2f_lw_axi_master_rvalid                                      : out std_logic;                                         -- rvalid
			hps_0_h2f_lw_axi_master_rready                                      : in  std_logic                      := 'X';             -- rready
			clk_0_clk_clk                                                       : in  std_logic                      := 'X';             -- clk
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			IN_DISPATCHER_clock_reset_reset_bridge_in_reset_reset               : in  std_logic                      := 'X';             -- reset
			IN_DISPATCHER_CSR_address                                           : out std_logic_vector(2 downto 0);                      -- address
			IN_DISPATCHER_CSR_write                                             : out std_logic;                                         -- write
			IN_DISPATCHER_CSR_read                                              : out std_logic;                                         -- read
			IN_DISPATCHER_CSR_readdata                                          : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			IN_DISPATCHER_CSR_writedata                                         : out std_logic_vector(31 downto 0);                     -- writedata
			IN_DISPATCHER_CSR_byteenable                                        : out std_logic_vector(3 downto 0);                      -- byteenable
			IN_DISPATCHER_Descriptor_Slave_write                                : out std_logic;                                         -- write
			IN_DISPATCHER_Descriptor_Slave_writedata                            : out std_logic_vector(127 downto 0);                    -- writedata
			IN_DISPATCHER_Descriptor_Slave_byteenable                           : out std_logic_vector(15 downto 0);                     -- byteenable
			IN_DISPATCHER_Descriptor_Slave_waitrequest                          : in  std_logic                      := 'X';             -- waitrequest
			QU_DISPATCHER_CSR_address                                           : out std_logic_vector(2 downto 0);                      -- address
			QU_DISPATCHER_CSR_write                                             : out std_logic;                                         -- write
			QU_DISPATCHER_CSR_read                                              : out std_logic;                                         -- read
			QU_DISPATCHER_CSR_readdata                                          : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			QU_DISPATCHER_CSR_writedata                                         : out std_logic_vector(31 downto 0);                     -- writedata
			QU_DISPATCHER_CSR_byteenable                                        : out std_logic_vector(3 downto 0);                      -- byteenable
			QU_DISPATCHER_Descriptor_Slave_write                                : out std_logic;                                         -- write
			QU_DISPATCHER_Descriptor_Slave_writedata                            : out std_logic_vector(127 downto 0);                    -- writedata
			QU_DISPATCHER_Descriptor_Slave_byteenable                           : out std_logic_vector(15 downto 0);                     -- byteenable
			QU_DISPATCHER_Descriptor_Slave_waitrequest                          : in  std_logic                      := 'X';             -- waitrequest
			recCtrl_0_recCtrlMM_write                                           : out std_logic;                                         -- write
			recCtrl_0_recCtrlMM_writedata                                       : out std_logic_vector(7 downto 0)                       -- writedata
		);
	end component soc_mm_interconnect_1;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal rfreceive_0_idatafifo_valid                                  : std_logic;                      -- RFReceive_0:rfRec_i_valid -> IN_DATA_FIFO:in_valid
	signal rfreceive_0_idatafifo_data                                   : std_logic_vector(15 downto 0);  -- RFReceive_0:rfRec_i_data -> IN_DATA_FIFO:in_data
	signal rfreceive_0_idatafifo_ready                                  : std_logic;                      -- IN_DATA_FIFO:in_ready -> RFReceive_0:rfRec_i_ready
	signal rfreceive_0_qdatafifo_valid                                  : std_logic;                      -- RFReceive_0:rfRec_q_valid -> QU_DATA_FIFO:in_valid
	signal rfreceive_0_qdatafifo_data                                   : std_logic_vector(15 downto 0);  -- RFReceive_0:rfRec_q_data -> QU_DATA_FIFO:in_data
	signal rfreceive_0_qdatafifo_ready                                  : std_logic;                      -- QU_DATA_FIFO:in_ready -> RFReceive_0:rfRec_q_ready
	signal in_write_master_response_source_valid                        : std_logic;                      -- IN_WRITE_MASTER:src_response_valid -> IN_DISPATCHER:snk_write_master_valid
	signal in_write_master_response_source_data                         : std_logic_vector(255 downto 0); -- IN_WRITE_MASTER:src_response_data -> IN_DISPATCHER:snk_write_master_data
	signal in_write_master_response_source_ready                        : std_logic;                      -- IN_DISPATCHER:snk_write_master_ready -> IN_WRITE_MASTER:src_response_ready
	signal qu_write_master_response_source_valid                        : std_logic;                      -- QU_WRITE_MASTER:src_response_valid -> QU_DISPATCHER:snk_write_master_valid
	signal qu_write_master_response_source_data                         : std_logic_vector(255 downto 0); -- QU_WRITE_MASTER:src_response_data -> QU_DISPATCHER:snk_write_master_data
	signal qu_write_master_response_source_ready                        : std_logic;                      -- QU_DISPATCHER:snk_write_master_ready -> QU_WRITE_MASTER:src_response_ready
	signal in_dispatcher_write_command_source_valid                     : std_logic;                      -- IN_DISPATCHER:src_write_master_valid -> IN_WRITE_MASTER:snk_command_valid
	signal in_dispatcher_write_command_source_data                      : std_logic_vector(255 downto 0); -- IN_DISPATCHER:src_write_master_data -> IN_WRITE_MASTER:snk_command_data
	signal in_dispatcher_write_command_source_ready                     : std_logic;                      -- IN_WRITE_MASTER:snk_command_ready -> IN_DISPATCHER:src_write_master_ready
	signal qu_dispatcher_write_command_source_valid                     : std_logic;                      -- QU_DISPATCHER:src_write_master_valid -> QU_WRITE_MASTER:snk_command_valid
	signal qu_dispatcher_write_command_source_data                      : std_logic_vector(255 downto 0); -- QU_DISPATCHER:src_write_master_data -> QU_WRITE_MASTER:snk_command_data
	signal qu_dispatcher_write_command_source_ready                     : std_logic;                      -- QU_WRITE_MASTER:snk_command_ready -> QU_DISPATCHER:src_write_master_ready
	signal in_data_fifo_out_valid                                       : std_logic;                      -- IN_DATA_FIFO:out_valid -> IN_WRITE_MASTER:snk_valid
	signal in_data_fifo_out_data                                        : std_logic_vector(15 downto 0);  -- IN_DATA_FIFO:out_data -> IN_WRITE_MASTER:snk_data
	signal in_data_fifo_out_ready                                       : std_logic;                      -- IN_WRITE_MASTER:snk_ready -> IN_DATA_FIFO:out_ready
	signal qu_data_fifo_out_valid                                       : std_logic;                      -- QU_DATA_FIFO:out_valid -> QU_WRITE_MASTER:snk_valid
	signal qu_data_fifo_out_data                                        : std_logic_vector(15 downto 0);  -- QU_DATA_FIFO:out_data -> QU_WRITE_MASTER:snk_data
	signal qu_data_fifo_out_ready                                       : std_logic;                      -- QU_WRITE_MASTER:snk_ready -> QU_DATA_FIFO:out_ready
	signal rfreceive_0_idatafifoclk_clk                                 : std_logic;                      -- RFReceive_0:rfRec_i_clk -> [IN_DATA_FIFO:in_clk, rst_controller:clk]
	signal rfreceive_0_qdatafifoclk_clk                                 : std_logic;                      -- RFReceive_0:rfRec_q_clk -> [QU_DATA_FIFO:in_clk, rst_controller_002:clk]
	signal in_write_master_data_write_master_waitrequest                : std_logic;                      -- mm_interconnect_0:IN_WRITE_MASTER_Data_Write_Master_waitrequest -> IN_WRITE_MASTER:master_waitrequest
	signal in_write_master_data_write_master_address                    : std_logic_vector(31 downto 0);  -- IN_WRITE_MASTER:master_address -> mm_interconnect_0:IN_WRITE_MASTER_Data_Write_Master_address
	signal in_write_master_data_write_master_byteenable                 : std_logic_vector(1 downto 0);   -- IN_WRITE_MASTER:master_byteenable -> mm_interconnect_0:IN_WRITE_MASTER_Data_Write_Master_byteenable
	signal in_write_master_data_write_master_write                      : std_logic;                      -- IN_WRITE_MASTER:master_write -> mm_interconnect_0:IN_WRITE_MASTER_Data_Write_Master_write
	signal in_write_master_data_write_master_writedata                  : std_logic_vector(15 downto 0);  -- IN_WRITE_MASTER:master_writedata -> mm_interconnect_0:IN_WRITE_MASTER_Data_Write_Master_writedata
	signal qu_write_master_data_write_master_waitrequest                : std_logic;                      -- mm_interconnect_0:QU_WRITE_MASTER_Data_Write_Master_waitrequest -> QU_WRITE_MASTER:master_waitrequest
	signal qu_write_master_data_write_master_address                    : std_logic_vector(31 downto 0);  -- QU_WRITE_MASTER:master_address -> mm_interconnect_0:QU_WRITE_MASTER_Data_Write_Master_address
	signal qu_write_master_data_write_master_byteenable                 : std_logic_vector(1 downto 0);   -- QU_WRITE_MASTER:master_byteenable -> mm_interconnect_0:QU_WRITE_MASTER_Data_Write_Master_byteenable
	signal qu_write_master_data_write_master_write                      : std_logic;                      -- QU_WRITE_MASTER:master_write -> mm_interconnect_0:QU_WRITE_MASTER_Data_Write_Master_write
	signal qu_write_master_data_write_master_writedata                  : std_logic_vector(15 downto 0);  -- QU_WRITE_MASTER:master_writedata -> mm_interconnect_0:QU_WRITE_MASTER_Data_Write_Master_writedata
	signal mm_interconnect_0_hps_0_f2h_sdram0_data_waitrequest          : std_logic;                      -- hps_0:f2h_sdram0_WAITREQUEST -> mm_interconnect_0:hps_0_f2h_sdram0_data_waitrequest
	signal mm_interconnect_0_hps_0_f2h_sdram0_data_address              : std_logic_vector(28 downto 0);  -- mm_interconnect_0:hps_0_f2h_sdram0_data_address -> hps_0:f2h_sdram0_ADDRESS
	signal mm_interconnect_0_hps_0_f2h_sdram0_data_byteenable           : std_logic_vector(7 downto 0);   -- mm_interconnect_0:hps_0_f2h_sdram0_data_byteenable -> hps_0:f2h_sdram0_BYTEENABLE
	signal mm_interconnect_0_hps_0_f2h_sdram0_data_write                : std_logic;                      -- mm_interconnect_0:hps_0_f2h_sdram0_data_write -> hps_0:f2h_sdram0_WRITE
	signal mm_interconnect_0_hps_0_f2h_sdram0_data_writedata            : std_logic_vector(63 downto 0);  -- mm_interconnect_0:hps_0_f2h_sdram0_data_writedata -> hps_0:f2h_sdram0_WRITEDATA
	signal mm_interconnect_0_hps_0_f2h_sdram0_data_burstcount           : std_logic_vector(7 downto 0);   -- mm_interconnect_0:hps_0_f2h_sdram0_data_burstcount -> hps_0:f2h_sdram0_BURSTCOUNT
	signal hps_0_h2f_lw_axi_master_awburst                              : std_logic_vector(1 downto 0);   -- hps_0:h2f_lw_AWBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awburst
	signal hps_0_h2f_lw_axi_master_arlen                                : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_ARLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlen
	signal hps_0_h2f_lw_axi_master_wstrb                                : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_WSTRB -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wstrb
	signal hps_0_h2f_lw_axi_master_wready                               : std_logic;                      -- mm_interconnect_1:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	signal hps_0_h2f_lw_axi_master_rid                                  : std_logic_vector(11 downto 0);  -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	signal hps_0_h2f_lw_axi_master_rready                               : std_logic;                      -- hps_0:h2f_lw_RREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_rready
	signal hps_0_h2f_lw_axi_master_awlen                                : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_AWLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlen
	signal hps_0_h2f_lw_axi_master_wid                                  : std_logic_vector(11 downto 0);  -- hps_0:h2f_lw_WID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wid
	signal hps_0_h2f_lw_axi_master_arcache                              : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_ARCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arcache
	signal hps_0_h2f_lw_axi_master_wvalid                               : std_logic;                      -- hps_0:h2f_lw_WVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wvalid
	signal hps_0_h2f_lw_axi_master_araddr                               : std_logic_vector(20 downto 0);  -- hps_0:h2f_lw_ARADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_araddr
	signal hps_0_h2f_lw_axi_master_arprot                               : std_logic_vector(2 downto 0);   -- hps_0:h2f_lw_ARPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arprot
	signal hps_0_h2f_lw_axi_master_awprot                               : std_logic_vector(2 downto 0);   -- hps_0:h2f_lw_AWPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awprot
	signal hps_0_h2f_lw_axi_master_wdata                                : std_logic_vector(31 downto 0);  -- hps_0:h2f_lw_WDATA -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wdata
	signal hps_0_h2f_lw_axi_master_arvalid                              : std_logic;                      -- hps_0:h2f_lw_ARVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arvalid
	signal hps_0_h2f_lw_axi_master_awcache                              : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_AWCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awcache
	signal hps_0_h2f_lw_axi_master_arid                                 : std_logic_vector(11 downto 0);  -- hps_0:h2f_lw_ARID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arid
	signal hps_0_h2f_lw_axi_master_arlock                               : std_logic_vector(1 downto 0);   -- hps_0:h2f_lw_ARLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlock
	signal hps_0_h2f_lw_axi_master_awlock                               : std_logic_vector(1 downto 0);   -- hps_0:h2f_lw_AWLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlock
	signal hps_0_h2f_lw_axi_master_awaddr                               : std_logic_vector(20 downto 0);  -- hps_0:h2f_lw_AWADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awaddr
	signal hps_0_h2f_lw_axi_master_bresp                                : std_logic_vector(1 downto 0);   -- mm_interconnect_1:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	signal hps_0_h2f_lw_axi_master_arready                              : std_logic;                      -- mm_interconnect_1:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	signal hps_0_h2f_lw_axi_master_rdata                                : std_logic_vector(31 downto 0);  -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	signal hps_0_h2f_lw_axi_master_awready                              : std_logic;                      -- mm_interconnect_1:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	signal hps_0_h2f_lw_axi_master_arburst                              : std_logic_vector(1 downto 0);   -- hps_0:h2f_lw_ARBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arburst
	signal hps_0_h2f_lw_axi_master_arsize                               : std_logic_vector(2 downto 0);   -- hps_0:h2f_lw_ARSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arsize
	signal hps_0_h2f_lw_axi_master_bready                               : std_logic;                      -- hps_0:h2f_lw_BREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_bready
	signal hps_0_h2f_lw_axi_master_rlast                                : std_logic;                      -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	signal hps_0_h2f_lw_axi_master_wlast                                : std_logic;                      -- hps_0:h2f_lw_WLAST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wlast
	signal hps_0_h2f_lw_axi_master_rresp                                : std_logic_vector(1 downto 0);   -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	signal hps_0_h2f_lw_axi_master_awid                                 : std_logic_vector(11 downto 0);  -- hps_0:h2f_lw_AWID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awid
	signal hps_0_h2f_lw_axi_master_bid                                  : std_logic_vector(11 downto 0);  -- mm_interconnect_1:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	signal hps_0_h2f_lw_axi_master_bvalid                               : std_logic;                      -- mm_interconnect_1:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	signal hps_0_h2f_lw_axi_master_awsize                               : std_logic_vector(2 downto 0);   -- hps_0:h2f_lw_AWSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awsize
	signal hps_0_h2f_lw_axi_master_awvalid                              : std_logic;                      -- hps_0:h2f_lw_AWVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awvalid
	signal hps_0_h2f_lw_axi_master_rvalid                               : std_logic;                      -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	signal mm_interconnect_1_in_dispatcher_csr_readdata                 : std_logic_vector(31 downto 0);  -- IN_DISPATCHER:csr_readdata -> mm_interconnect_1:IN_DISPATCHER_CSR_readdata
	signal mm_interconnect_1_in_dispatcher_csr_address                  : std_logic_vector(2 downto 0);   -- mm_interconnect_1:IN_DISPATCHER_CSR_address -> IN_DISPATCHER:csr_address
	signal mm_interconnect_1_in_dispatcher_csr_read                     : std_logic;                      -- mm_interconnect_1:IN_DISPATCHER_CSR_read -> IN_DISPATCHER:csr_read
	signal mm_interconnect_1_in_dispatcher_csr_byteenable               : std_logic_vector(3 downto 0);   -- mm_interconnect_1:IN_DISPATCHER_CSR_byteenable -> IN_DISPATCHER:csr_byteenable
	signal mm_interconnect_1_in_dispatcher_csr_write                    : std_logic;                      -- mm_interconnect_1:IN_DISPATCHER_CSR_write -> IN_DISPATCHER:csr_write
	signal mm_interconnect_1_in_dispatcher_csr_writedata                : std_logic_vector(31 downto 0);  -- mm_interconnect_1:IN_DISPATCHER_CSR_writedata -> IN_DISPATCHER:csr_writedata
	signal mm_interconnect_1_qu_dispatcher_csr_readdata                 : std_logic_vector(31 downto 0);  -- QU_DISPATCHER:csr_readdata -> mm_interconnect_1:QU_DISPATCHER_CSR_readdata
	signal mm_interconnect_1_qu_dispatcher_csr_address                  : std_logic_vector(2 downto 0);   -- mm_interconnect_1:QU_DISPATCHER_CSR_address -> QU_DISPATCHER:csr_address
	signal mm_interconnect_1_qu_dispatcher_csr_read                     : std_logic;                      -- mm_interconnect_1:QU_DISPATCHER_CSR_read -> QU_DISPATCHER:csr_read
	signal mm_interconnect_1_qu_dispatcher_csr_byteenable               : std_logic_vector(3 downto 0);   -- mm_interconnect_1:QU_DISPATCHER_CSR_byteenable -> QU_DISPATCHER:csr_byteenable
	signal mm_interconnect_1_qu_dispatcher_csr_write                    : std_logic;                      -- mm_interconnect_1:QU_DISPATCHER_CSR_write -> QU_DISPATCHER:csr_write
	signal mm_interconnect_1_qu_dispatcher_csr_writedata                : std_logic_vector(31 downto 0);  -- mm_interconnect_1:QU_DISPATCHER_CSR_writedata -> QU_DISPATCHER:csr_writedata
	signal mm_interconnect_1_in_dispatcher_descriptor_slave_waitrequest : std_logic;                      -- IN_DISPATCHER:descriptor_waitrequest -> mm_interconnect_1:IN_DISPATCHER_Descriptor_Slave_waitrequest
	signal mm_interconnect_1_in_dispatcher_descriptor_slave_byteenable  : std_logic_vector(15 downto 0);  -- mm_interconnect_1:IN_DISPATCHER_Descriptor_Slave_byteenable -> IN_DISPATCHER:descriptor_byteenable
	signal mm_interconnect_1_in_dispatcher_descriptor_slave_write       : std_logic;                      -- mm_interconnect_1:IN_DISPATCHER_Descriptor_Slave_write -> IN_DISPATCHER:descriptor_write
	signal mm_interconnect_1_in_dispatcher_descriptor_slave_writedata   : std_logic_vector(127 downto 0); -- mm_interconnect_1:IN_DISPATCHER_Descriptor_Slave_writedata -> IN_DISPATCHER:descriptor_writedata
	signal mm_interconnect_1_qu_dispatcher_descriptor_slave_waitrequest : std_logic;                      -- QU_DISPATCHER:descriptor_waitrequest -> mm_interconnect_1:QU_DISPATCHER_Descriptor_Slave_waitrequest
	signal mm_interconnect_1_qu_dispatcher_descriptor_slave_byteenable  : std_logic_vector(15 downto 0);  -- mm_interconnect_1:QU_DISPATCHER_Descriptor_Slave_byteenable -> QU_DISPATCHER:descriptor_byteenable
	signal mm_interconnect_1_qu_dispatcher_descriptor_slave_write       : std_logic;                      -- mm_interconnect_1:QU_DISPATCHER_Descriptor_Slave_write -> QU_DISPATCHER:descriptor_write
	signal mm_interconnect_1_qu_dispatcher_descriptor_slave_writedata   : std_logic_vector(127 downto 0); -- mm_interconnect_1:QU_DISPATCHER_Descriptor_Slave_writedata -> QU_DISPATCHER:descriptor_writedata
	signal mm_interconnect_1_recctrl_0_recctrlmm_write                  : std_logic;                      -- mm_interconnect_1:recCtrl_0_recCtrlMM_write -> recCtrl_0:write_en
	signal mm_interconnect_1_recctrl_0_recctrlmm_writedata              : std_logic_vector(7 downto 0);   -- mm_interconnect_1:recCtrl_0_recCtrlMM_writedata -> recCtrl_0:write_data
	signal rst_controller_reset_out_reset                               : std_logic;                      -- rst_controller:reset_out -> rst_controller_reset_out_reset:in
	signal rst_controller_001_reset_out_reset                           : std_logic;                      -- rst_controller_001:reset_out -> [IN_DISPATCHER:reset, IN_WRITE_MASTER:reset, QU_DISPATCHER:reset, QU_WRITE_MASTER:reset, RFReceive_0:reset, mm_interconnect_0:IN_WRITE_MASTER_Clock_reset_reset_bridge_in_reset_reset, mm_interconnect_1:IN_DISPATCHER_clock_reset_reset_bridge_in_reset_reset, recCtrl_0:reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_002_reset_out_reset                           : std_logic;                      -- rst_controller_002:reset_out -> rst_controller_002_reset_out_reset:in
	signal rst_controller_003_reset_out_reset                           : std_logic;                      -- rst_controller_003:reset_out -> [mm_interconnect_0:hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]
	signal hps_0_h2f_reset_reset                                        : std_logic;                      -- hps_0:h2f_rst_n -> hps_0_h2f_reset_reset:in
	signal reset_reset_n_ports_inv                                      : std_logic;                      -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal rst_controller_reset_out_reset_ports_inv                     : std_logic;                      -- rst_controller_reset_out_reset:inv -> IN_DATA_FIFO:in_reset_n
	signal rst_controller_001_reset_out_reset_ports_inv                 : std_logic;                      -- rst_controller_001_reset_out_reset:inv -> [IN_DATA_FIFO:out_reset_n, QU_DATA_FIFO:out_reset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                 : std_logic;                      -- rst_controller_002_reset_out_reset:inv -> QU_DATA_FIFO:in_reset_n
	signal hps_0_h2f_reset_reset_ports_inv                              : std_logic;                      -- hps_0_h2f_reset_reset:inv -> rst_controller_003:reset_in0

begin

	in_data_fifo : component altera_avalon_dc_fifo
		generic map (
			SYMBOLS_PER_BEAT   => 2,
			BITS_PER_SYMBOL    => 8,
			FIFO_DEPTH         => 2048,
			CHANNEL_WIDTH      => 0,
			ERROR_WIDTH        => 0,
			USE_PACKETS        => 0,
			USE_IN_FILL_LEVEL  => 0,
			USE_OUT_FILL_LEVEL => 0,
			WR_SYNC_DEPTH      => 16,
			RD_SYNC_DEPTH      => 16
		)
		port map (
			in_clk            => rfreceive_0_idatafifoclk_clk,                 --        in_clk.clk
			in_reset_n        => rst_controller_reset_out_reset_ports_inv,     --  in_clk_reset.reset_n
			out_clk           => clk_clk,                                      --       out_clk.clk
			out_reset_n       => rst_controller_001_reset_out_reset_ports_inv, -- out_clk_reset.reset_n
			in_data           => rfreceive_0_idatafifo_data,                   --            in.data
			in_valid          => rfreceive_0_idatafifo_valid,                  --              .valid
			in_ready          => rfreceive_0_idatafifo_ready,                  --              .ready
			out_data          => in_data_fifo_out_data,                        --           out.data
			out_valid         => in_data_fifo_out_valid,                       --              .valid
			out_ready         => in_data_fifo_out_ready,                       --              .ready
			in_csr_address    => '0',                                          --   (terminated)
			in_csr_read       => '0',                                          --   (terminated)
			in_csr_write      => '0',                                          --   (terminated)
			in_csr_readdata   => open,                                         --   (terminated)
			in_csr_writedata  => "00000000000000000000000000000000",           --   (terminated)
			out_csr_address   => '0',                                          --   (terminated)
			out_csr_read      => '0',                                          --   (terminated)
			out_csr_write     => '0',                                          --   (terminated)
			out_csr_readdata  => open,                                         --   (terminated)
			out_csr_writedata => "00000000000000000000000000000000",           --   (terminated)
			in_startofpacket  => '0',                                          --   (terminated)
			in_endofpacket    => '0',                                          --   (terminated)
			out_startofpacket => open,                                         --   (terminated)
			out_endofpacket   => open                                          --   (terminated)
		);

	in_dispatcher : component dispatcher
		generic map (
			MODE                        => 2,
			RESPONSE_PORT               => 2,
			DESCRIPTOR_FIFO_DEPTH       => 8,
			ENHANCED_FEATURES           => 0,
			DESCRIPTOR_WIDTH            => 128,
			DESCRIPTOR_BYTEENABLE_WIDTH => 16
		)
		port map (
			clk                     => clk_clk,                                                                                                                                                                                                                                                            --                clock.clk
			reset                   => rst_controller_001_reset_out_reset,                                                                                                                                                                                                                                 --          clock_reset.reset
			csr_writedata           => mm_interconnect_1_in_dispatcher_csr_writedata,                                                                                                                                                                                                                      --                  CSR.writedata
			csr_write               => mm_interconnect_1_in_dispatcher_csr_write,                                                                                                                                                                                                                          --                     .write
			csr_byteenable          => mm_interconnect_1_in_dispatcher_csr_byteenable,                                                                                                                                                                                                                     --                     .byteenable
			csr_readdata            => mm_interconnect_1_in_dispatcher_csr_readdata,                                                                                                                                                                                                                       --                     .readdata
			csr_read                => mm_interconnect_1_in_dispatcher_csr_read,                                                                                                                                                                                                                           --                     .read
			csr_address             => mm_interconnect_1_in_dispatcher_csr_address,                                                                                                                                                                                                                        --                     .address
			descriptor_write        => mm_interconnect_1_in_dispatcher_descriptor_slave_write,                                                                                                                                                                                                             --     Descriptor_Slave.write
			descriptor_waitrequest  => mm_interconnect_1_in_dispatcher_descriptor_slave_waitrequest,                                                                                                                                                                                                       --                     .waitrequest
			descriptor_writedata    => mm_interconnect_1_in_dispatcher_descriptor_slave_writedata,                                                                                                                                                                                                         --                     .writedata
			descriptor_byteenable   => mm_interconnect_1_in_dispatcher_descriptor_slave_byteenable,                                                                                                                                                                                                        --                     .byteenable
			src_write_master_data   => in_dispatcher_write_command_source_data,                                                                                                                                                                                                                            -- Write_Command_Source.data
			src_write_master_valid  => in_dispatcher_write_command_source_valid,                                                                                                                                                                                                                           --                     .valid
			src_write_master_ready  => in_dispatcher_write_command_source_ready,                                                                                                                                                                                                                           --                     .ready
			snk_write_master_data   => in_write_master_response_source_data,                                                                                                                                                                                                                               --  Write_Response_Sink.data
			snk_write_master_valid  => in_write_master_response_source_valid,                                                                                                                                                                                                                              --                     .valid
			snk_write_master_ready  => in_write_master_response_source_ready,                                                                                                                                                                                                                              --                     .ready
			csr_irq                 => open,                                                                                                                                                                                                                                                               --              csr_irq.irq
			src_response_data       => open,                                                                                                                                                                                                                                                               --          (terminated)
			src_response_valid      => open,                                                                                                                                                                                                                                                               --          (terminated)
			src_response_ready      => '0',                                                                                                                                                                                                                                                                --          (terminated)
			mm_response_waitrequest => open,                                                                                                                                                                                                                                                               --          (terminated)
			mm_response_byteenable  => "0000",                                                                                                                                                                                                                                                             --          (terminated)
			mm_response_address     => '0',                                                                                                                                                                                                                                                                --          (terminated)
			mm_response_readdata    => open,                                                                                                                                                                                                                                                               --          (terminated)
			mm_response_read        => '0',                                                                                                                                                                                                                                                                --          (terminated)
			src_read_master_data    => open,                                                                                                                                                                                                                                                               --          (terminated)
			src_read_master_valid   => open,                                                                                                                                                                                                                                                               --          (terminated)
			src_read_master_ready   => '0',                                                                                                                                                                                                                                                                --          (terminated)
			snk_read_master_data    => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --          (terminated)
			snk_read_master_valid   => '0',                                                                                                                                                                                                                                                                --          (terminated)
			snk_read_master_ready   => open                                                                                                                                                                                                                                                                --          (terminated)
		);

	in_write_master : component write_master
		generic map (
			DATA_WIDTH                     => 16,
			LENGTH_WIDTH                   => 32,
			FIFO_DEPTH                     => 128,
			STRIDE_ENABLE                  => 0,
			BURST_ENABLE                   => 0,
			PACKET_ENABLE                  => 0,
			ERROR_ENABLE                   => 0,
			ERROR_WIDTH                    => 8,
			BYTE_ENABLE_WIDTH              => 2,
			BYTE_ENABLE_WIDTH_LOG2         => 1,
			ADDRESS_WIDTH                  => 32,
			FIFO_DEPTH_LOG2                => 7,
			SYMBOL_WIDTH                   => 8,
			NUMBER_OF_SYMBOLS              => 2,
			NUMBER_OF_SYMBOLS_LOG2         => 1,
			MAX_BURST_COUNT_WIDTH          => 1,
			UNALIGNED_ACCESSES_ENABLE      => 0,
			ONLY_FULL_ACCESS_ENABLE        => 0,
			BURST_WRAPPING_SUPPORT         => 0,
			PROGRAMMABLE_BURST_ENABLE      => 0,
			MAX_BURST_COUNT                => 1,
			FIFO_SPEED_OPTIMIZATION        => 1,
			STRIDE_WIDTH                   => 1,
			ACTUAL_BYTES_TRANSFERRED_WIDTH => 32
		)
		port map (
			clk                => clk_clk,                                       --             Clock.clk
			reset              => rst_controller_001_reset_out_reset,            --       Clock_reset.reset
			master_address     => in_write_master_data_write_master_address,     -- Data_Write_Master.address
			master_write       => in_write_master_data_write_master_write,       --                  .write
			master_byteenable  => in_write_master_data_write_master_byteenable,  --                  .byteenable
			master_writedata   => in_write_master_data_write_master_writedata,   --                  .writedata
			master_waitrequest => in_write_master_data_write_master_waitrequest, --                  .waitrequest
			snk_data           => in_data_fifo_out_data,                         --         Data_Sink.data
			snk_valid          => in_data_fifo_out_valid,                        --                  .valid
			snk_ready          => in_data_fifo_out_ready,                        --                  .ready
			snk_command_data   => in_dispatcher_write_command_source_data,       --      Command_Sink.data
			snk_command_valid  => in_dispatcher_write_command_source_valid,      --                  .valid
			snk_command_ready  => in_dispatcher_write_command_source_ready,      --                  .ready
			src_response_data  => in_write_master_response_source_data,          --   Response_Source.data
			src_response_valid => in_write_master_response_source_valid,         --                  .valid
			src_response_ready => in_write_master_response_source_ready,         --                  .ready
			master_burstcount  => open,                                          --       (terminated)
			snk_sop            => '0',                                           --       (terminated)
			snk_eop            => '0',                                           --       (terminated)
			snk_empty          => '0',                                           --       (terminated)
			snk_error          => "00000000"                                     --       (terminated)
		);

	qu_data_fifo : component altera_avalon_dc_fifo
		generic map (
			SYMBOLS_PER_BEAT   => 2,
			BITS_PER_SYMBOL    => 8,
			FIFO_DEPTH         => 2048,
			CHANNEL_WIDTH      => 0,
			ERROR_WIDTH        => 0,
			USE_PACKETS        => 0,
			USE_IN_FILL_LEVEL  => 0,
			USE_OUT_FILL_LEVEL => 0,
			WR_SYNC_DEPTH      => 16,
			RD_SYNC_DEPTH      => 16
		)
		port map (
			in_clk            => rfreceive_0_qdatafifoclk_clk,                 --        in_clk.clk
			in_reset_n        => rst_controller_002_reset_out_reset_ports_inv, --  in_clk_reset.reset_n
			out_clk           => clk_clk,                                      --       out_clk.clk
			out_reset_n       => rst_controller_001_reset_out_reset_ports_inv, -- out_clk_reset.reset_n
			in_data           => rfreceive_0_qdatafifo_data,                   --            in.data
			in_valid          => rfreceive_0_qdatafifo_valid,                  --              .valid
			in_ready          => rfreceive_0_qdatafifo_ready,                  --              .ready
			out_data          => qu_data_fifo_out_data,                        --           out.data
			out_valid         => qu_data_fifo_out_valid,                       --              .valid
			out_ready         => qu_data_fifo_out_ready,                       --              .ready
			in_csr_address    => '0',                                          --   (terminated)
			in_csr_read       => '0',                                          --   (terminated)
			in_csr_write      => '0',                                          --   (terminated)
			in_csr_readdata   => open,                                         --   (terminated)
			in_csr_writedata  => "00000000000000000000000000000000",           --   (terminated)
			out_csr_address   => '0',                                          --   (terminated)
			out_csr_read      => '0',                                          --   (terminated)
			out_csr_write     => '0',                                          --   (terminated)
			out_csr_readdata  => open,                                         --   (terminated)
			out_csr_writedata => "00000000000000000000000000000000",           --   (terminated)
			in_startofpacket  => '0',                                          --   (terminated)
			in_endofpacket    => '0',                                          --   (terminated)
			out_startofpacket => open,                                         --   (terminated)
			out_endofpacket   => open                                          --   (terminated)
		);

	qu_dispatcher : component dispatcher
		generic map (
			MODE                        => 2,
			RESPONSE_PORT               => 2,
			DESCRIPTOR_FIFO_DEPTH       => 8,
			ENHANCED_FEATURES           => 0,
			DESCRIPTOR_WIDTH            => 128,
			DESCRIPTOR_BYTEENABLE_WIDTH => 16
		)
		port map (
			clk                     => clk_clk,                                                                                                                                                                                                                                                            --                clock.clk
			reset                   => rst_controller_001_reset_out_reset,                                                                                                                                                                                                                                 --          clock_reset.reset
			csr_writedata           => mm_interconnect_1_qu_dispatcher_csr_writedata,                                                                                                                                                                                                                      --                  CSR.writedata
			csr_write               => mm_interconnect_1_qu_dispatcher_csr_write,                                                                                                                                                                                                                          --                     .write
			csr_byteenable          => mm_interconnect_1_qu_dispatcher_csr_byteenable,                                                                                                                                                                                                                     --                     .byteenable
			csr_readdata            => mm_interconnect_1_qu_dispatcher_csr_readdata,                                                                                                                                                                                                                       --                     .readdata
			csr_read                => mm_interconnect_1_qu_dispatcher_csr_read,                                                                                                                                                                                                                           --                     .read
			csr_address             => mm_interconnect_1_qu_dispatcher_csr_address,                                                                                                                                                                                                                        --                     .address
			descriptor_write        => mm_interconnect_1_qu_dispatcher_descriptor_slave_write,                                                                                                                                                                                                             --     Descriptor_Slave.write
			descriptor_waitrequest  => mm_interconnect_1_qu_dispatcher_descriptor_slave_waitrequest,                                                                                                                                                                                                       --                     .waitrequest
			descriptor_writedata    => mm_interconnect_1_qu_dispatcher_descriptor_slave_writedata,                                                                                                                                                                                                         --                     .writedata
			descriptor_byteenable   => mm_interconnect_1_qu_dispatcher_descriptor_slave_byteenable,                                                                                                                                                                                                        --                     .byteenable
			src_write_master_data   => qu_dispatcher_write_command_source_data,                                                                                                                                                                                                                            -- Write_Command_Source.data
			src_write_master_valid  => qu_dispatcher_write_command_source_valid,                                                                                                                                                                                                                           --                     .valid
			src_write_master_ready  => qu_dispatcher_write_command_source_ready,                                                                                                                                                                                                                           --                     .ready
			snk_write_master_data   => qu_write_master_response_source_data,                                                                                                                                                                                                                               --  Write_Response_Sink.data
			snk_write_master_valid  => qu_write_master_response_source_valid,                                                                                                                                                                                                                              --                     .valid
			snk_write_master_ready  => qu_write_master_response_source_ready,                                                                                                                                                                                                                              --                     .ready
			csr_irq                 => open,                                                                                                                                                                                                                                                               --              csr_irq.irq
			src_response_data       => open,                                                                                                                                                                                                                                                               --          (terminated)
			src_response_valid      => open,                                                                                                                                                                                                                                                               --          (terminated)
			src_response_ready      => '0',                                                                                                                                                                                                                                                                --          (terminated)
			mm_response_waitrequest => open,                                                                                                                                                                                                                                                               --          (terminated)
			mm_response_byteenable  => "0000",                                                                                                                                                                                                                                                             --          (terminated)
			mm_response_address     => '0',                                                                                                                                                                                                                                                                --          (terminated)
			mm_response_readdata    => open,                                                                                                                                                                                                                                                               --          (terminated)
			mm_response_read        => '0',                                                                                                                                                                                                                                                                --          (terminated)
			src_read_master_data    => open,                                                                                                                                                                                                                                                               --          (terminated)
			src_read_master_valid   => open,                                                                                                                                                                                                                                                               --          (terminated)
			src_read_master_ready   => '0',                                                                                                                                                                                                                                                                --          (terminated)
			snk_read_master_data    => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --          (terminated)
			snk_read_master_valid   => '0',                                                                                                                                                                                                                                                                --          (terminated)
			snk_read_master_ready   => open                                                                                                                                                                                                                                                                --          (terminated)
		);

	qu_write_master : component write_master
		generic map (
			DATA_WIDTH                     => 16,
			LENGTH_WIDTH                   => 32,
			FIFO_DEPTH                     => 128,
			STRIDE_ENABLE                  => 0,
			BURST_ENABLE                   => 0,
			PACKET_ENABLE                  => 0,
			ERROR_ENABLE                   => 0,
			ERROR_WIDTH                    => 8,
			BYTE_ENABLE_WIDTH              => 2,
			BYTE_ENABLE_WIDTH_LOG2         => 1,
			ADDRESS_WIDTH                  => 32,
			FIFO_DEPTH_LOG2                => 7,
			SYMBOL_WIDTH                   => 8,
			NUMBER_OF_SYMBOLS              => 2,
			NUMBER_OF_SYMBOLS_LOG2         => 1,
			MAX_BURST_COUNT_WIDTH          => 1,
			UNALIGNED_ACCESSES_ENABLE      => 0,
			ONLY_FULL_ACCESS_ENABLE        => 0,
			BURST_WRAPPING_SUPPORT         => 0,
			PROGRAMMABLE_BURST_ENABLE      => 0,
			MAX_BURST_COUNT                => 1,
			FIFO_SPEED_OPTIMIZATION        => 1,
			STRIDE_WIDTH                   => 1,
			ACTUAL_BYTES_TRANSFERRED_WIDTH => 32
		)
		port map (
			clk                => clk_clk,                                       --             Clock.clk
			reset              => rst_controller_001_reset_out_reset,            --       Clock_reset.reset
			master_address     => qu_write_master_data_write_master_address,     -- Data_Write_Master.address
			master_write       => qu_write_master_data_write_master_write,       --                  .write
			master_byteenable  => qu_write_master_data_write_master_byteenable,  --                  .byteenable
			master_writedata   => qu_write_master_data_write_master_writedata,   --                  .writedata
			master_waitrequest => qu_write_master_data_write_master_waitrequest, --                  .waitrequest
			snk_data           => qu_data_fifo_out_data,                         --         Data_Sink.data
			snk_valid          => qu_data_fifo_out_valid,                        --                  .valid
			snk_ready          => qu_data_fifo_out_ready,                        --                  .ready
			snk_command_data   => qu_dispatcher_write_command_source_data,       --      Command_Sink.data
			snk_command_valid  => qu_dispatcher_write_command_source_valid,      --                  .valid
			snk_command_ready  => qu_dispatcher_write_command_source_ready,      --                  .ready
			src_response_data  => qu_write_master_response_source_data,          --   Response_Source.data
			src_response_valid => qu_write_master_response_source_valid,         --                  .valid
			src_response_ready => qu_write_master_response_source_ready,         --                  .ready
			master_burstcount  => open,                                          --       (terminated)
			snk_sop            => '0',                                           --       (terminated)
			snk_eop            => '0',                                           --       (terminated)
			snk_empty          => '0',                                           --       (terminated)
			snk_error          => "00000000"                                     --       (terminated)
		);

	rfreceive_0 : component RFReceive
		port map (
			clk           => clk_clk,                            --        clock.clk
			reset         => rst_controller_001_reset_out_reset, --        reset.reset
			RXCLK         => rfrec_rxclock,                      --      conduit.rxclock
			RXD           => rfrec_rxdata,                       --             .rxdata
			RXEN          => rfrec_rxenable,                     --             .rxenable
			RXIQSEL       => rfrec_rxiq,                         --             .rxiq
			RecEnable     => rfrec_recen,                        --             .recen
			LED           => rfrec_testled,                      --             .testled
			rfRec_i_data  => rfreceive_0_idatafifo_data,         --    IDataFIFO.data
			rfRec_i_ready => rfreceive_0_idatafifo_ready,        --             .ready
			rfRec_i_valid => rfreceive_0_idatafifo_valid,        --             .valid
			rfRec_q_data  => rfreceive_0_qdatafifo_data,         --    QDataFIFO.data
			rfRec_q_ready => rfreceive_0_qdatafifo_ready,        --             .ready
			rfRec_q_valid => rfreceive_0_qdatafifo_valid,        --             .valid
			rfRec_i_clk   => rfreceive_0_idatafifoclk_clk,       -- IDataFIFOCLK.clk
			rfRec_q_clk   => rfreceive_0_qdatafifoclk_clk        -- QDataFIFOCLK.clk
		);

	hps_0 : component soc_hps_0
		generic map (
			F2S_Width => 0,
			S2F_Width => 0
		)
		port map (
			mem_a                  => memory_mem_a,                                        --            memory.mem_a
			mem_ba                 => memory_mem_ba,                                       --                  .mem_ba
			mem_ck                 => memory_mem_ck,                                       --                  .mem_ck
			mem_ck_n               => memory_mem_ck_n,                                     --                  .mem_ck_n
			mem_cke                => memory_mem_cke,                                      --                  .mem_cke
			mem_cs_n               => memory_mem_cs_n,                                     --                  .mem_cs_n
			mem_ras_n              => memory_mem_ras_n,                                    --                  .mem_ras_n
			mem_cas_n              => memory_mem_cas_n,                                    --                  .mem_cas_n
			mem_we_n               => memory_mem_we_n,                                     --                  .mem_we_n
			mem_reset_n            => memory_mem_reset_n,                                  --                  .mem_reset_n
			mem_dq                 => memory_mem_dq,                                       --                  .mem_dq
			mem_dqs                => memory_mem_dqs,                                      --                  .mem_dqs
			mem_dqs_n              => memory_mem_dqs_n,                                    --                  .mem_dqs_n
			mem_odt                => memory_mem_odt,                                      --                  .mem_odt
			mem_dm                 => memory_mem_dm,                                       --                  .mem_dm
			oct_rzqin              => memory_oct_rzqin,                                    --                  .oct_rzqin
			h2f_rst_n              => hps_0_h2f_reset_reset,                               --         h2f_reset.reset_n
			f2h_sdram0_clk         => clk_clk,                                             --  f2h_sdram0_clock.clk
			f2h_sdram0_ADDRESS     => mm_interconnect_0_hps_0_f2h_sdram0_data_address,     --   f2h_sdram0_data.address
			f2h_sdram0_BURSTCOUNT  => mm_interconnect_0_hps_0_f2h_sdram0_data_burstcount,  --                  .burstcount
			f2h_sdram0_WAITREQUEST => mm_interconnect_0_hps_0_f2h_sdram0_data_waitrequest, --                  .waitrequest
			f2h_sdram0_WRITEDATA   => mm_interconnect_0_hps_0_f2h_sdram0_data_writedata,   --                  .writedata
			f2h_sdram0_BYTEENABLE  => mm_interconnect_0_hps_0_f2h_sdram0_data_byteenable,  --                  .byteenable
			f2h_sdram0_WRITE       => mm_interconnect_0_hps_0_f2h_sdram0_data_write,       --                  .write
			h2f_lw_axi_clk         => clk_clk,                                             --  h2f_lw_axi_clock.clk
			h2f_lw_AWID            => hps_0_h2f_lw_axi_master_awid,                        -- h2f_lw_axi_master.awid
			h2f_lw_AWADDR          => hps_0_h2f_lw_axi_master_awaddr,                      --                  .awaddr
			h2f_lw_AWLEN           => hps_0_h2f_lw_axi_master_awlen,                       --                  .awlen
			h2f_lw_AWSIZE          => hps_0_h2f_lw_axi_master_awsize,                      --                  .awsize
			h2f_lw_AWBURST         => hps_0_h2f_lw_axi_master_awburst,                     --                  .awburst
			h2f_lw_AWLOCK          => hps_0_h2f_lw_axi_master_awlock,                      --                  .awlock
			h2f_lw_AWCACHE         => hps_0_h2f_lw_axi_master_awcache,                     --                  .awcache
			h2f_lw_AWPROT          => hps_0_h2f_lw_axi_master_awprot,                      --                  .awprot
			h2f_lw_AWVALID         => hps_0_h2f_lw_axi_master_awvalid,                     --                  .awvalid
			h2f_lw_AWREADY         => hps_0_h2f_lw_axi_master_awready,                     --                  .awready
			h2f_lw_WID             => hps_0_h2f_lw_axi_master_wid,                         --                  .wid
			h2f_lw_WDATA           => hps_0_h2f_lw_axi_master_wdata,                       --                  .wdata
			h2f_lw_WSTRB           => hps_0_h2f_lw_axi_master_wstrb,                       --                  .wstrb
			h2f_lw_WLAST           => hps_0_h2f_lw_axi_master_wlast,                       --                  .wlast
			h2f_lw_WVALID          => hps_0_h2f_lw_axi_master_wvalid,                      --                  .wvalid
			h2f_lw_WREADY          => hps_0_h2f_lw_axi_master_wready,                      --                  .wready
			h2f_lw_BID             => hps_0_h2f_lw_axi_master_bid,                         --                  .bid
			h2f_lw_BRESP           => hps_0_h2f_lw_axi_master_bresp,                       --                  .bresp
			h2f_lw_BVALID          => hps_0_h2f_lw_axi_master_bvalid,                      --                  .bvalid
			h2f_lw_BREADY          => hps_0_h2f_lw_axi_master_bready,                      --                  .bready
			h2f_lw_ARID            => hps_0_h2f_lw_axi_master_arid,                        --                  .arid
			h2f_lw_ARADDR          => hps_0_h2f_lw_axi_master_araddr,                      --                  .araddr
			h2f_lw_ARLEN           => hps_0_h2f_lw_axi_master_arlen,                       --                  .arlen
			h2f_lw_ARSIZE          => hps_0_h2f_lw_axi_master_arsize,                      --                  .arsize
			h2f_lw_ARBURST         => hps_0_h2f_lw_axi_master_arburst,                     --                  .arburst
			h2f_lw_ARLOCK          => hps_0_h2f_lw_axi_master_arlock,                      --                  .arlock
			h2f_lw_ARCACHE         => hps_0_h2f_lw_axi_master_arcache,                     --                  .arcache
			h2f_lw_ARPROT          => hps_0_h2f_lw_axi_master_arprot,                      --                  .arprot
			h2f_lw_ARVALID         => hps_0_h2f_lw_axi_master_arvalid,                     --                  .arvalid
			h2f_lw_ARREADY         => hps_0_h2f_lw_axi_master_arready,                     --                  .arready
			h2f_lw_RID             => hps_0_h2f_lw_axi_master_rid,                         --                  .rid
			h2f_lw_RDATA           => hps_0_h2f_lw_axi_master_rdata,                       --                  .rdata
			h2f_lw_RRESP           => hps_0_h2f_lw_axi_master_rresp,                       --                  .rresp
			h2f_lw_RLAST           => hps_0_h2f_lw_axi_master_rlast,                       --                  .rlast
			h2f_lw_RVALID          => hps_0_h2f_lw_axi_master_rvalid,                      --                  .rvalid
			h2f_lw_RREADY          => hps_0_h2f_lw_axi_master_rready                       --                  .rready
		);

	recctrl_0 : component recCtrl
		port map (
			clk        => clk_clk,                                         --     clock.clk
			reset      => rst_controller_001_reset_out_reset,              --     reset.reset
			RecEnable  => reccontrol_enrec,                                --   conduit.enrec
			write_data => mm_interconnect_1_recctrl_0_recctrlmm_writedata, -- recCtrlMM.writedata
			write_en   => mm_interconnect_1_recctrl_0_recctrlmm_write      --          .write
		);

	mm_interconnect_0 : component soc_mm_interconnect_0
		port map (
			clk_0_clk_clk                                                      => clk_clk,                                             --                                                    clk_0_clk.clk
			hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset => rst_controller_003_reset_out_reset,                  -- hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset.reset
			IN_WRITE_MASTER_Clock_reset_reset_bridge_in_reset_reset            => rst_controller_001_reset_out_reset,                  --            IN_WRITE_MASTER_Clock_reset_reset_bridge_in_reset.reset
			IN_WRITE_MASTER_Data_Write_Master_address                          => in_write_master_data_write_master_address,           --                            IN_WRITE_MASTER_Data_Write_Master.address
			IN_WRITE_MASTER_Data_Write_Master_waitrequest                      => in_write_master_data_write_master_waitrequest,       --                                                             .waitrequest
			IN_WRITE_MASTER_Data_Write_Master_byteenable                       => in_write_master_data_write_master_byteenable,        --                                                             .byteenable
			IN_WRITE_MASTER_Data_Write_Master_write                            => in_write_master_data_write_master_write,             --                                                             .write
			IN_WRITE_MASTER_Data_Write_Master_writedata                        => in_write_master_data_write_master_writedata,         --                                                             .writedata
			QU_WRITE_MASTER_Data_Write_Master_address                          => qu_write_master_data_write_master_address,           --                            QU_WRITE_MASTER_Data_Write_Master.address
			QU_WRITE_MASTER_Data_Write_Master_waitrequest                      => qu_write_master_data_write_master_waitrequest,       --                                                             .waitrequest
			QU_WRITE_MASTER_Data_Write_Master_byteenable                       => qu_write_master_data_write_master_byteenable,        --                                                             .byteenable
			QU_WRITE_MASTER_Data_Write_Master_write                            => qu_write_master_data_write_master_write,             --                                                             .write
			QU_WRITE_MASTER_Data_Write_Master_writedata                        => qu_write_master_data_write_master_writedata,         --                                                             .writedata
			hps_0_f2h_sdram0_data_address                                      => mm_interconnect_0_hps_0_f2h_sdram0_data_address,     --                                        hps_0_f2h_sdram0_data.address
			hps_0_f2h_sdram0_data_write                                        => mm_interconnect_0_hps_0_f2h_sdram0_data_write,       --                                                             .write
			hps_0_f2h_sdram0_data_writedata                                    => mm_interconnect_0_hps_0_f2h_sdram0_data_writedata,   --                                                             .writedata
			hps_0_f2h_sdram0_data_burstcount                                   => mm_interconnect_0_hps_0_f2h_sdram0_data_burstcount,  --                                                             .burstcount
			hps_0_f2h_sdram0_data_byteenable                                   => mm_interconnect_0_hps_0_f2h_sdram0_data_byteenable,  --                                                             .byteenable
			hps_0_f2h_sdram0_data_waitrequest                                  => mm_interconnect_0_hps_0_f2h_sdram0_data_waitrequest  --                                                             .waitrequest
		);

	mm_interconnect_1 : component soc_mm_interconnect_1
		port map (
			hps_0_h2f_lw_axi_master_awid                                        => hps_0_h2f_lw_axi_master_awid,                                 --                                       hps_0_h2f_lw_axi_master.awid
			hps_0_h2f_lw_axi_master_awaddr                                      => hps_0_h2f_lw_axi_master_awaddr,                               --                                                              .awaddr
			hps_0_h2f_lw_axi_master_awlen                                       => hps_0_h2f_lw_axi_master_awlen,                                --                                                              .awlen
			hps_0_h2f_lw_axi_master_awsize                                      => hps_0_h2f_lw_axi_master_awsize,                               --                                                              .awsize
			hps_0_h2f_lw_axi_master_awburst                                     => hps_0_h2f_lw_axi_master_awburst,                              --                                                              .awburst
			hps_0_h2f_lw_axi_master_awlock                                      => hps_0_h2f_lw_axi_master_awlock,                               --                                                              .awlock
			hps_0_h2f_lw_axi_master_awcache                                     => hps_0_h2f_lw_axi_master_awcache,                              --                                                              .awcache
			hps_0_h2f_lw_axi_master_awprot                                      => hps_0_h2f_lw_axi_master_awprot,                               --                                                              .awprot
			hps_0_h2f_lw_axi_master_awvalid                                     => hps_0_h2f_lw_axi_master_awvalid,                              --                                                              .awvalid
			hps_0_h2f_lw_axi_master_awready                                     => hps_0_h2f_lw_axi_master_awready,                              --                                                              .awready
			hps_0_h2f_lw_axi_master_wid                                         => hps_0_h2f_lw_axi_master_wid,                                  --                                                              .wid
			hps_0_h2f_lw_axi_master_wdata                                       => hps_0_h2f_lw_axi_master_wdata,                                --                                                              .wdata
			hps_0_h2f_lw_axi_master_wstrb                                       => hps_0_h2f_lw_axi_master_wstrb,                                --                                                              .wstrb
			hps_0_h2f_lw_axi_master_wlast                                       => hps_0_h2f_lw_axi_master_wlast,                                --                                                              .wlast
			hps_0_h2f_lw_axi_master_wvalid                                      => hps_0_h2f_lw_axi_master_wvalid,                               --                                                              .wvalid
			hps_0_h2f_lw_axi_master_wready                                      => hps_0_h2f_lw_axi_master_wready,                               --                                                              .wready
			hps_0_h2f_lw_axi_master_bid                                         => hps_0_h2f_lw_axi_master_bid,                                  --                                                              .bid
			hps_0_h2f_lw_axi_master_bresp                                       => hps_0_h2f_lw_axi_master_bresp,                                --                                                              .bresp
			hps_0_h2f_lw_axi_master_bvalid                                      => hps_0_h2f_lw_axi_master_bvalid,                               --                                                              .bvalid
			hps_0_h2f_lw_axi_master_bready                                      => hps_0_h2f_lw_axi_master_bready,                               --                                                              .bready
			hps_0_h2f_lw_axi_master_arid                                        => hps_0_h2f_lw_axi_master_arid,                                 --                                                              .arid
			hps_0_h2f_lw_axi_master_araddr                                      => hps_0_h2f_lw_axi_master_araddr,                               --                                                              .araddr
			hps_0_h2f_lw_axi_master_arlen                                       => hps_0_h2f_lw_axi_master_arlen,                                --                                                              .arlen
			hps_0_h2f_lw_axi_master_arsize                                      => hps_0_h2f_lw_axi_master_arsize,                               --                                                              .arsize
			hps_0_h2f_lw_axi_master_arburst                                     => hps_0_h2f_lw_axi_master_arburst,                              --                                                              .arburst
			hps_0_h2f_lw_axi_master_arlock                                      => hps_0_h2f_lw_axi_master_arlock,                               --                                                              .arlock
			hps_0_h2f_lw_axi_master_arcache                                     => hps_0_h2f_lw_axi_master_arcache,                              --                                                              .arcache
			hps_0_h2f_lw_axi_master_arprot                                      => hps_0_h2f_lw_axi_master_arprot,                               --                                                              .arprot
			hps_0_h2f_lw_axi_master_arvalid                                     => hps_0_h2f_lw_axi_master_arvalid,                              --                                                              .arvalid
			hps_0_h2f_lw_axi_master_arready                                     => hps_0_h2f_lw_axi_master_arready,                              --                                                              .arready
			hps_0_h2f_lw_axi_master_rid                                         => hps_0_h2f_lw_axi_master_rid,                                  --                                                              .rid
			hps_0_h2f_lw_axi_master_rdata                                       => hps_0_h2f_lw_axi_master_rdata,                                --                                                              .rdata
			hps_0_h2f_lw_axi_master_rresp                                       => hps_0_h2f_lw_axi_master_rresp,                                --                                                              .rresp
			hps_0_h2f_lw_axi_master_rlast                                       => hps_0_h2f_lw_axi_master_rlast,                                --                                                              .rlast
			hps_0_h2f_lw_axi_master_rvalid                                      => hps_0_h2f_lw_axi_master_rvalid,                               --                                                              .rvalid
			hps_0_h2f_lw_axi_master_rready                                      => hps_0_h2f_lw_axi_master_rready,                               --                                                              .rready
			clk_0_clk_clk                                                       => clk_clk,                                                      --                                                     clk_0_clk.clk
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_003_reset_out_reset,                           -- hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			IN_DISPATCHER_clock_reset_reset_bridge_in_reset_reset               => rst_controller_001_reset_out_reset,                           --               IN_DISPATCHER_clock_reset_reset_bridge_in_reset.reset
			IN_DISPATCHER_CSR_address                                           => mm_interconnect_1_in_dispatcher_csr_address,                  --                                             IN_DISPATCHER_CSR.address
			IN_DISPATCHER_CSR_write                                             => mm_interconnect_1_in_dispatcher_csr_write,                    --                                                              .write
			IN_DISPATCHER_CSR_read                                              => mm_interconnect_1_in_dispatcher_csr_read,                     --                                                              .read
			IN_DISPATCHER_CSR_readdata                                          => mm_interconnect_1_in_dispatcher_csr_readdata,                 --                                                              .readdata
			IN_DISPATCHER_CSR_writedata                                         => mm_interconnect_1_in_dispatcher_csr_writedata,                --                                                              .writedata
			IN_DISPATCHER_CSR_byteenable                                        => mm_interconnect_1_in_dispatcher_csr_byteenable,               --                                                              .byteenable
			IN_DISPATCHER_Descriptor_Slave_write                                => mm_interconnect_1_in_dispatcher_descriptor_slave_write,       --                                IN_DISPATCHER_Descriptor_Slave.write
			IN_DISPATCHER_Descriptor_Slave_writedata                            => mm_interconnect_1_in_dispatcher_descriptor_slave_writedata,   --                                                              .writedata
			IN_DISPATCHER_Descriptor_Slave_byteenable                           => mm_interconnect_1_in_dispatcher_descriptor_slave_byteenable,  --                                                              .byteenable
			IN_DISPATCHER_Descriptor_Slave_waitrequest                          => mm_interconnect_1_in_dispatcher_descriptor_slave_waitrequest, --                                                              .waitrequest
			QU_DISPATCHER_CSR_address                                           => mm_interconnect_1_qu_dispatcher_csr_address,                  --                                             QU_DISPATCHER_CSR.address
			QU_DISPATCHER_CSR_write                                             => mm_interconnect_1_qu_dispatcher_csr_write,                    --                                                              .write
			QU_DISPATCHER_CSR_read                                              => mm_interconnect_1_qu_dispatcher_csr_read,                     --                                                              .read
			QU_DISPATCHER_CSR_readdata                                          => mm_interconnect_1_qu_dispatcher_csr_readdata,                 --                                                              .readdata
			QU_DISPATCHER_CSR_writedata                                         => mm_interconnect_1_qu_dispatcher_csr_writedata,                --                                                              .writedata
			QU_DISPATCHER_CSR_byteenable                                        => mm_interconnect_1_qu_dispatcher_csr_byteenable,               --                                                              .byteenable
			QU_DISPATCHER_Descriptor_Slave_write                                => mm_interconnect_1_qu_dispatcher_descriptor_slave_write,       --                                QU_DISPATCHER_Descriptor_Slave.write
			QU_DISPATCHER_Descriptor_Slave_writedata                            => mm_interconnect_1_qu_dispatcher_descriptor_slave_writedata,   --                                                              .writedata
			QU_DISPATCHER_Descriptor_Slave_byteenable                           => mm_interconnect_1_qu_dispatcher_descriptor_slave_byteenable,  --                                                              .byteenable
			QU_DISPATCHER_Descriptor_Slave_waitrequest                          => mm_interconnect_1_qu_dispatcher_descriptor_slave_waitrequest, --                                                              .waitrequest
			recCtrl_0_recCtrlMM_write                                           => mm_interconnect_1_recctrl_0_recctrlmm_write,                  --                                           recCtrl_0_recCtrlMM.write
			recCtrl_0_recCtrlMM_writedata                                       => mm_interconnect_1_recctrl_0_recctrlmm_writedata               --                                                              .writedata
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => rfreceive_0_idatafifoclk_clk,   --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => rfreceive_0_qdatafifoclk_clk,       --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_003 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_0_h2f_reset_reset_ports_inv,    -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

	hps_0_h2f_reset_reset_ports_inv <= not hps_0_h2f_reset_reset;

end architecture rtl; -- of soc
